`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
nBWkdC6e7Fy2AHsDMMYIwua19I/8ampGCVKfZKZEEquvGcK/QthUPmcNsTHSRiDeRNAY7QpqoAjI
Y00/IgD+Dw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eFOXXSZHhC72U7yv9eXEqPTFD5mKDeM/flBAkXGqEbTLwBpL4uFm4lc7ujktgt9kJG3iA2Jo0uL/
VlAI4gNy+T+8hFpiCGw5KEhy9Vc9fzoGJEIbYWlYSKabVx6usZDKOdJJgOFhgpysRlnzmMnRKK1F
gWIGRenSxsfpilXa5QI=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
S+dVFBludpj6IonNToIKx+WZsCy5cjeuHZJyTUb9LJu08jba7BK9sEpu+SOJ4hoxyzZmVMFP4nnA
Rn74joUR6lZgmqcam8r5MIyA2vYqpgNwNYAN6RXrGHdoIHU1QR/HNxOP6y8gk2dENkv/OJsMYY5/
sgGwnSESY6PfUkFWLhDt5rbAeqKQi6eIk2HL/MSgwdE8zn4ILombREeYxZHRw0VB9K+SjbLWOFpY
Z8FNBSj5FF0VHRcwqtcyP56a77O33LxQQR1EfGSg6nWnb0GN77XUMyjqW7dreFiOle1bL2FDPq8R
IlTit2jl1AGyujoxdvlt8GSnnScDmysbDeJR/w==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OYWZfcLYfEA9xtB1o5+F1vR8vP5fbJ1t1v9l1yWh+LLbgndznCn40HLA/5mP+iZ0ugmjeHI95IUh
GqAnAU7/74RzIiF9PbasPClDpHeZGsF+XNCoMwzREBy4np9VmD/PVHdbFaZwwYi17/+tGeyqQJ3/
DNhbyVj2zIzE0aPUuPLsCYhky8e4jiryqNichx52F28eTPppHfSODhoZiwgTWxpxaQ8SZUvkyvRd
wHGKgOj7pO9iUZemfFda31LfRG7+9AjVA2oal72pdsSmHMDZi9BMXar8ZfdJhxqwEBi6nn2S6cYA
xvazbYYgTxGv88/1AXVSf8fvz2Pxd/Zwj4BuGA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OOHITo+qPQ+AuOSufWzolP1KTlC0iDKCyIUPZUBdtoU74OIjItPVd8Q2Iw2pMK9qRcaYPS8oK1TB
R0KPhsClrukMOSnuCq1Tm9h8VSjXD0HZtVfN5tVNHU+e9gISv9NCFAwWD+BLgD2QxftXfgq/c7YG
wQdlInV+aXf9sIfzg1cQA1WtR7LYrEaui9X9asPxLx1M5aVM5rjCOPPJrsMukZ42uxE1pu5abVoT
jzF8eQqsu9sXTeYd/UgGOvXzYUblU65REeddRKOpr/FJqe+4i7WK+eSIQpI60GqZsKzRCiDTwPi/
HuwO8ix4vxwtUTGm2aN6Z5+IfKTlT0OOWjzRSg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TDK5yH4x6uFYmGzDvYc5q2U7AxGad3Mw1+yuQxjr7QeR93LeYRfmPRyhIV/unNJAnaKAzI/0sURH
Dzg0ILuuiGRb+a/U3xDljetdpQsAWHi1esC7JXwO1i+hMX8bdyflwSvmj6iZ1OBIB0VnhlxH4kti
HggJnuEGbV4T2yTmSkw=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RQn2qn8HlwJ+JfEQn4eLFBGllaDnvPclcK7vvB/J4wmRM+y89+x9XUNCzVWvXUXHpeeOSz1VkItT
om+bK8KKS8dzVaDDLkqw+XbeiJ43wJ0Yf/m0PR8D12CBqAVrXERYQr6+jDCiDWdCR/OdpS0B1LnQ
F+uAvHLJJtTcSi5Z0o4J6+JA+mCIghFN22fgfy5S4XBDHkskeUW18FAroctUdANFYvwomFNUum7F
EiDzbzt2mCp+W/gX0Z97jvwJ+C47oVT6IY9vgSjZ9HhipfVB00D9qgWAEJYnlmnxvQC2Wt3BCMdO
PL86p0nfdrsinX1bT4Z5pAzVUB5CjLhww69nYw==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LDCPTyLEkGzmRP98uXGsg/a+VW9cQm7UhDCD0/9tWJF7OHI+u/OIF8y2Ar0jrKBioRg2oWRVUwXW
LqAQEoGfVc2VIaCdlvGLGrKP9Dah1ZgjYaK27BWn6UMpOoURG3d0LuYTsr2JFZ93rxRWLHt7MPXn
8fw2irSXEXpxZvOSZ+0eQURb1o5ww7vja7U1grE5wwM97t6aoKma1Nmj/O0jnwJLHSSqUAdX5ski
J16fWynYraD8HxUJwWMOctqEvkM+lDn521JhjNLNuVPfE+oQVjlWtJpzKoc2ko+Or5Qp9hfgCBZP
N/58VOcPYG2XCw/xY+E+tbPtU6lOSp4i/6wYcg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 133696)
`protect data_block
WWJrYdvC04a1lVZGHN2w9er3u+GOyDXdqpJClDuKN4vJBR8X8lKe0qJGTN62PfB/4ZlH1OVFpRaQ
I+XAA5/eu9SEUm7n1OhaHPI65GmTU5qd3lbmogvf19RN0LQoES3HbskWPDeNi59OgaiWcKcGCmNg
OpqTwP5lbmTt1a2hJ9mP+0QPSRA72U565qe3vC+/Pp9hOY5SMjExkcDxWz1ZIFXNLnJqp1rYQOa3
HAyJB3i4j3l8n9LMXNQABaxLgUGqs/ycJe9KwUImaRDouTBc+gH3ANlvTcWhxNvYwyU608nwyBrU
JgFBAmIdqbGgGEuUxmwg+D7bJLPBQ56WwSs3Jo+X4HpeUaQLkuE3VRRq9RV7rauoD9CbTw7nXF02
D7GEGazFW20ePP9U6biyYTtw6XSEFGORMBOuD3EV7e2RSXBlkrXlLEmDatmMvxboHYvbGhAN1zss
RuPKDvVUPaClw++8Bb2Nqny73BN0v/NIpm7MfA3Y8VRG2aZToVpYZ0fH53mSIRCoMp79HD8WZZWC
I2yjf92VqAcHLBtHFsGTVjTQ/0Tb9Kn7MdVyQYflgkIr8mZyzMFyBbq7qMqetJI+jN/l5GiFKIx/
rcNpoHs+twyMThwDFVvHHu8cT9XuuKFTTL7rknzWWkEc7YxdDnMFiyvmxXm4nL6NAvAkcAnfm++X
7vmS5lK8K1zt2bTlCo4NsUAXX8mpE4CWhHvfN5YsESUChOfjKIVwTR9Zu3jQBTYJGOncFnjM9hyh
3OQF2E573FLBYbqU6eGkJ0yMvAFcf6ZNGSEoLGHISKCG8RUYwyUznrGmkTVGsKwCorfYSYKhgVOx
hUaMXxj3EcMMeuNG3txl5yxGUbQY/bJyTiighrptfcaRE4RJzywwwS3VjTKdI6olshkcio5AJiGS
IKVhgIjKjGKlhSApiw9FfRcMqR8xpsFK/bUIgnfgT6rSeK742UiM9K7XNLuzxtTthrTTJuMIYpFJ
0PzzVYO6fu1Bhq2UoRrgSB+oymKgE1Lx1p/KMFBemsPCkwJaiMH2oTW0fhTnW4HsQPUdVd/GZdpf
7uOfxbbX+CdqOFDT1VaiIQvXG7S1tL0UnVYqbkg0ORdpqWw7SOp9JeElA9jnytFVvAHjjrzJxYeN
54XwHhkPAoZpHwNp2cT2EdVT/rghnNReLQ03q+nIP2L0Ld6vQILAMAmttRJLFbud/aniE2Yg2CnH
T0L9tmV8JYuDsHR9QEt0Q78OzwzHuN0QKjT59UEVHaKBeZVzigQ5ULXfPCuqNEbm+KF/Gq38SLpD
0GQlF9x5x9UI1/jefWi1qJCY0IrXawa3m5VZ+qjQJEQVIu0Dr113wmPYN3lsAi0cKon+hV3WkNFe
G9K/prNC9lNPRhcy1b7SexlvVvEn61vu5QGU6KgW18ZMg+ENWBCHQ2s/gy1XJ5+ZymQQrhHYEt82
glrwv7pcmazztdZJlj2HDcvHu/etCf8a7fkY80VW0qQX1Y1AcK0/GNYDkA6nogdN1N42tvdQrTfD
KU24Rem5VDUpf8paiojtYk4SflAGbOilxb9GJy+NDdAuB3UDiNOK1nc8oNgGc2r/gZ48sl6AVa8E
HTx3MKqJSpsCb6r6Oi7t9HcFkM5ACctU2nknkCrjwgzJnVYEcHAKGB7bhOF1MjzePDYsKhJyTITq
iOM2PRClfPv+Kh93RygZ6EJYI3wfacqMG1/oLZ7PSQuBYFBCHnESBHQ1FJvq5MwwPnSCHbgXwirz
w9O5X4u7cg0JbC/CDNLTNIgUgJ7OYNbmThTrJNEHP7LfvGwOF48p+zWLL8+54xO6zkx5glEeF907
Ofb/WX6cdBVn/4P1YI33kiiD5X6OrliWTz100ebXyDduPqhbFqYIX8jgnZqjKbi8to8EKulSaVGn
qHPbt/Z9Bcr6CCMBaaZQj+CQu0LCDhbbWGcwwuN2pQSAqWD0E8aY5EfTgQiJbXuPLSSfzify6EDm
CZIB96JYM9lzzfXQ33ofr9mkXu3ZZgHpUMEEPgOkSJifCfGBhHLzdS9WzH3Hl9d9LMKnBIVs4Yle
j8IuNj0DIPJjAhRctaUbCHvX2wJq3Wu0+Zz+v+h2YM3HZSeDvsLPsl2HXOzZXURX1wh6V4xQCZMW
S+Hdz7cTNYcmHW1E6gC9RK44RD8F7EfECa8mNhEpIn2/bisdbDGmYtDRHIwLoB7rgUy9si2hFb+U
Ckyla8azoohiuT3CmegdPrRX5QNJbQL7VfE7ZdR8nW6vvfHQ95w1lqDBiNmRlIV90FPD4yuGThrX
7YGdvpiJLUiuxMk632WEK5T+D9IqSKfqEF5uzvJBuiEDhV4kjTzjHHzxr78uOIZpSprxBkTd6SF8
/637tPMWrZkx+Q81SNkko7OInFUUScjeGbpV/tfzzTZwcCK+xPv3CM4GVF2H9boVzZRis7yTr9IA
2Eaun/esXEKIMaSiL3NSuy1uc0aTdIFdFVDbzEm54XAO5jjyqmaTX3Yq4jfW2b6ndRJ9M9ku3VKU
+kM42Scs7gQq80XwLcL4bcP2BJnvS7BJIl8ANiSgSOAmQL6+99ZosLqzMTSr9s/dbNpZzZap1etK
bZMpQHgdupz0xITRgu9G7yY7aPl9oB34025AGjQe9JCDKMvXr6asbevQyfp7KB3A4soyyJ8LSnVS
4280U9sGJCw/UDkyMCBHyl1bqX6KDMb9tBtke1NhCGxoz0QUir4YEe1vyOaxG10uuIwvb1wxzwgf
Bivow74nLovUBbNgt/DfM2djwT864QuNFZFCmoVgW2emSFo7vmL7GDiJ6m8jJvY0nLpkpK7LFhL8
NiODmUXdFWb+PMt1vocAv5+w73SZHivwdb5QpMWpYbe7LYOFbrh6Wsj2tkjZMtDeSYgooiENiqes
QDXJzbg4ypyL7gYW+rEklYTMnUGB585KvnXdgdZtY8u3oHHf0jQZ+zQhqkztnPnRDM/4Cu++e2MS
TUSAcv1H/GoLiu+ouaoSOqPH+VJ01/aC6+O4/J1vR8zPky8bHJpk/yFNJin1Gw/5ZI01Q6Dms8zM
Hgbtf6B1GTvnmSGPafPe1YaMt52fv8iPRx0EhnsFEjXbUnb+cj99o3yRdu0M9ZMOPx5doErlicTT
ukXDb+BZV63zkTdAelMW2E+QlZTMGqkO2GzBAuXnJCPxuCq8Hc520z32Q0yc6ggENnUHRUEXwhO5
Ke7/UUHYW/rqFYvmvXKvhldYSCoLn02N/yFQErYC5jlDnddHzFmjQY9wWUEHSCPEzTiYOAoAx/ys
OGrZMEZ82W71p8AXB8z0jwUBgCLgC0QRx3VfLaTNGueryPZNgu9b6u3W5zqPHIN2pqVBDcBEPOLh
7Ahd1vtBKhr5PeJ9FefeEM698SvqMtSE3Xzlc97KNXj8BDJFAcPQmqlp+ic2TRw/MAextP/yg2tW
+vCnjAcq54i0DRJj/mwTydlQICC9UjRMLYBF8ogUKKhsGMlgMnioPXCzfuEirNedrmUuWohA3gRh
oUDfgK/x5/WqllTv2+4Ur6kFIei4SRbfhdxZ5Fs+yYM6ECQcVFkwR4YWJdKXQAqBn4yATWiy1bky
zepAttT6uVSwoJBwozzvmgLEAooUZy9dV+IkcLyH1ec2MRsi+gipSE3kitcCfUinODCRYq7T5dNY
xxrCH8nddbpsW7Jo+rC9Jo1th0tl3BpjqGqNjMyvuLdngEwk+uRsS//u22PfQkGxZizw/42RlShM
FqZWlsmbWf2w1jFTVhqf2onAMtpW5EzOZ5Oox6n3LcKqbt6gXKgjLOKj/f1quXJViLj2qk8ATcmi
YYqL9IfAB2ya6yt5TtYIlam11TK8bQTHB1RpNFamT+urTv7CGl4PIjioy+7xCSY3IMQKOyu85MD0
JQ2DmGi6g2Z4GCjeQAU6kNWcWprjhU/FRPaqvDeD1UhyqHO0tLm5q9kMQ834+DoqGWRa8oUYiDD6
K5btPu9N64nmnElBZeGXres4fHJ1sIzUWj8VVZcac4cviofxAdHVhK5jWpu1SJL8SxOxG92R/xiu
Edej21oMMNjYId8EzbnvpaajX1Em9GHUc7/lbjWVMDUE3juE7p2uq089Ulgx7K/T80x+HGm4l3wl
nM/EYDTdFxelyRsp9qUVqzlV2XCz76TdDoxSX3JEEZeZ0kgLDzpPKtAjN6cc1Zb1SonOx73TFdpc
9eO5zyJW6ld5T9zvs2J+qGeZAAJx+/zTLEvWyySVvWzibI8l+WKBh9eof6irdi4M9Jsw7ruDFZVz
w66/090bgfxT/JGc71PrWs4dhLikwZSF1AvcfvpS3UR/nzUeJyA33SHYn5FFoIDxGCvE+oeErebU
IRs9yLw95vcJgKB3HyabJi+1QnnqcDmuUixdgeZXNB+adHlH5elRJAgeOnHhF2MhTvK7mgS90WcE
lBoqUBD9JC2MVPDV/iBm0Lf/my6Bm9ckMLaxdbsPviZ6Bc94y8jqnTHFwQ+O3mrmFZwEh6As+J1h
DJs9vAlJ2d40ohqnADD2JUB+4Uek8swTcjCq2Oay5qLwjVTLWufPIDlpxy8JE1CTLaMGdcS9cWg0
6ZD0QkpWIK1fuhmTF6a1y7WaQDPiftMTRBBnpuIIkw0wekR4edgtYpxwKxPBrmqf1T+VY3oRl+u0
Tiy+3s6xCsh+DvjBngrpuRP6wrWxQKesOx8iD3UIm0myVh9G3IATQEu6vR0KAKkiy5VV3gUVVo2w
24/3JfOGOZ5uEC4GOGok3BUEM8vgneGT7ln5PMplBwVjq/1H7B4H7P571aXoKH59eaTy2EYlyJpk
RUD3LwMB6bz5C6TdEEZXodvQjb0WGXwNTcZ6VAttQm7FyeQ0NSQLzwkLdECbpp1rvLOoqMnXCnvK
4GrbXcEHTKyu6j+QrZx9gLmnUHySDNX9y4XCJu6eOCxN+bpFyV7OJq+T7ZUdrV56QQhrAT9f7O8x
Z9PgPmGNYABvhfYhBi8Ty1IQSUATC1WOe2I8ETga47jX/51rGH+PWKNfkDTCA0tzCPFv0OoM6jm+
Ih5qWXurCKH45CFOilvFDpUjuj/upsFJU0a9GvFeYuUME1kzWzBb0bNqDXsXqi7X6x+COE7R4axp
8TuYvPC4JWqREPu4iAtUqwWn6V5wYcUNB8uLJBi8qGEIl1T0k1ci74RHUfVKtYNV0bLb4OReFnJK
izoXMbloPp4jkcTBezEtip9JOpR4nhGnXPd6zfzT1NSpcvRa/5yB5lnsa541FPtS4TBhesGNoNau
7vFD0L96bqz2Q1o8fBTDqKFodbNi6++Moy3r7zdVQFcL7PG7EL9LQtkM8nVUnCPvGotVktv5/cX0
HbWslZI2h9TjBuHARKJmbda6kKauD56kz4QKes0ypjgElNoWZCNAnz6vt2Rk1ucCQBVEROBJHaJN
FWMZvVzMmVWA7Riv5m7kNV1Sfhuo5Xww+vYrAVRxDJ48fxFAXdP5OdFGA/2Du0inp+euZz/OovT+
YH8TkV3LZ+S1BCMDSuw6QUrZGDfAX3NeFnT8slHnzk9Eb1+M22t08E8ZxN7GS3diV2V4YsJTt9+I
97Ea350Q74SrY7EMYF7MjWZGobvo3wubNoD0gOuFa4ssqv9hBHI+gIUl9tyr+zXjIln6ypa5sRP3
Irk0fL3xhucbrNJuAjK11wLr+XFv7jY5bCut5n6aSqqmxC7bC+p2uKk+bV5G6Rb4o+ZQeTn6UPBB
lUoj17EMXDXeW3d3A8OGr/NX3buAcYkowp4TkVi7sgMCqZo3foFkCzfXDGkB45ji6PV4PLQRasMi
pWHqYCjYO67LjTHLVwGXp+4qSJ46IPlB/RTFRydmx+s+Ug2L0B+uAMX830kDo0mvBbS+Td313JHq
nYMQwdMXWA59uePiMIfbDSlFwbahDmg6UGsp8/UC90x8zW6CNYO4/854qOxZ2k28LO2HuVjs3hqJ
cKOWmwHwBzAPRY2/TzYVeDXmV+yru96Bx4JwoS09bFaGWjhjjE/HsiQAeHN59NGmBknDuAAmT3jk
A/VIele09Bdyn7CkSG45XcSoQAi6f6M/HcTmR5rDJZolZWe8RxU9nwHI35GQ0+C3B9MOpa1vwXNf
o+UKnWVwVCKKqOO1raY1wqgd/+tQONSamRheHlADqEFbRsvL8iz2cAer1JF8gSBGjbmLkOSRG/HV
39id1wzHmZz+VTERRpLyusN5o1ALFL83K/4NaryyhHs0E9TpvmJbg7hlTKh+45qJGMgeEIdV6Xdn
SizaRsT8ot9UnSBHik9l45dI11MjGI78DBSPtHHf5e4y+tol4HlGJLhYmBy3RDxj2l9thX8UUu+d
lrQP6CuLWvOGrCmTcKlFTdWGY4RTuzRJer6ibCiI5hjoDKB14tDYDOQ7wO29uQsgpEqB77f78qlD
U6TCE5vGT7o1bES3MuIlEFvv2hbOMagwFf7Ifu0MhOrwN33ba6P2RU5CJdzw4S4jwAKKqOQ/jUEz
1mD0kgV/YWdblnCAu2U3l8j7DVUP6n0I75Y4kEJkihQwO3WwiWnyzuHJvMQBhhKJOu18GZXic6Mg
U1JwjqhN603rA65fR4oqveIq/fcPlQbieO+U/LanBPtw+I94mWTgr0bN2XKh9zwr4TE+/lUzNZ2v
bSBFNUeErJT+flTyJLy7Jb5oJU8yTm/yTPqeZLO4qUwvlimAPC1RG6USrmc9aOiN/QK/WdnOJkwi
los33o9Wy3Hk9mrKLyxoaZETmG4sVVw/OJtWxuhJ4jRsN/Cg7Jf8/phRXe0B/6hvD/j378tBhdsC
wt7kR/w2MBKkQ/xHm+MInH37JGXJvG1WtO5SBRCoStOWHwlGRuO5fSnvY2V44c06yJCwLMna55vS
Y5HW2nhKh66QwRwC3cjOsVF4Or7NeeRBDl22xXHHW+c0F3zySB2ztTuATpu27bPAp/lISZ+262vt
HO05t82ukDEPt7vq5vO/YJyue8i5qaSxBBvZJvV5zkPtt8r0xXkqUsAdEktYJzwM+3PjTZXT36iW
MweZqhvrdEkSfaLuBDaVAUgpA+sFTWlYlgQnxwjoguA9hURdBgcRheSCYoC997GXiksco42dpYZN
a4tj/bwkvLStjFr5H9/u8EXPNDFQvrypPiiwny0dEEF1m3V+BJsMqXURhrmsrVR8rzwaLp4UfAHD
S3Etjt7BWZymSI85E+E5bn1/wIb+daJCpjbGZU+O/R9sfJsE7E1p/Af2DrdooJPx5FoKHXWPfCDs
Fi1Q8FSKf6cyw79WPB3mPEcI/xe8vGycYZMx49CBavwmxQV21Po7y3uR3BFH+KrNBnBBD0Rvf9R3
LxWYj+CYFH4y0e48wI2ogLF1f5n+eiPT6EkoB0mKQfZ/REumfGeDA/JprsKaHtis6Q3KJSmvk4y+
4V6bRG/H+9TW3nXo01GEEG4st0AhRg8mqLdXBl4V4uKD2nrScKs5YHpoFQFLJ0LSarw9pA0GIVUc
GfieUjgJO9M4crzE5KFZFbnFhTEeCF9onQ/zkG263QvReIfWBotSwjCTklHBG2n8QkwfGORBhPd+
9iwdnQZFfHcQhWbzWm1OsQwaZjQfAfndguDXXY4O1/jZ7AptaU8oLuSmTbfBjCBt9OjM2jojsqmH
IWqEkrYvJZSDDNG9dwp9rO6GAwRBw8zISfXmQF+BOFE/5UE1iHAm3G9n22R5xwhiNG/I3v4k3jHu
eMZfOBfQyD/2YP9GtPrRheyQVdUC0gidET5CeQFUlK5PH0u64s2H9C7XTM3YcE7oSW9Mt5Ac8qt/
JXsno36u3r9nTzv6IjMkoQtRsXgTByOOwJU+4vApYt1+4bF4NNZqwSgCrjaOzEjPaU3gY62bI+SR
dZUWRHLmcG8C6FmeglTzeSKDEe1NK13PdDCY2+O2h3V/0Om+ktb/IGGD+S0uvagnBykb3cXE1sOE
vnSV1Z4lnSbQ5x6pBFCM8fSOSAsRKy2vvAYhaSt7sOkfvU0aKQ2IQ2MVAyNMCnRdnYl2hoMsOJpE
D79eLP83PUF4srCQ4y5S5DJop+GtTzvdGJp3A+kZP7FqdDKTrRjlUXdfnRuQuaLdzDOfVy86M7hV
WoyuTmVvIUwF3xRWMOmEMioLG6+PLOHJMFd8mVBB1VWhuLoc5mBzjGMFQ7Tck99DCduDTNMowbea
RAWUVAzuF4jDfi+LKH1cvUGU7d7avg9p4+adOqoYoLu6CP28XMPf8KzsRS4H2YhMJGtnRscjMBZ5
enu9FhFpyvkpoklz5VLOB2guNHRZY7P3CA+fh1hp6jxWEVcUopzZo/kpJepoXlT2NA80e5h/+6IS
wbhYZpUTjxNRrjsuK2YUbvssxQhy8xDm2R8Eqpwo/Cys+kmbz0afBWjQWL7U7rdZyccEiyO5oOj9
8BfGNofV7Z4V1duu+7cnrNeMKmTRbRVdvCJuDFARxVwqdyfStci99nWHhjAhUz+Caf//2C9SiWvs
2GrX/+nbHgx/smeFM69jEYyx8FmVQPVPIPv0aNzg3ziHvdJnipZRAV7RqWT2nYFtdil+KFgNffW2
atoYZrOQlJJ1gS4CFwhYojuiF/ol0LECGnaSrk53ZkLPiPy7yjnfPO4ZRHF+LpZdlFqE511jyizB
u5bScIqgCkd3eVG2iLjqlwM+KVZmoiDCWKoN3duMsN2S3sFarTar4wCMA5NdRZoc36xmTi8hgRct
968E8+7YoOGaaUAiOZ++hH1OBsapVwo907vYJcNQD27HQMm4lwF9Lu+QBRBoUw82RMIyELNSXlI7
J9TKDEc8SYyAAErs4Z0ABo+m1WNyuNl4AtzkAg4FSK0CWEHQXq2QHgzCHpXPaJ0XnvaJynwZ6Pb3
Aov9rDK5jpNjUkoZxl6tHoa83YzOGZdUMJC22M8nosBSzY1SY0VdCvndfSpJ0fDwllv75WfoHgjM
VDmWbm35a9pvU0xeeciMwumaNljjx793FWqlFJ+vjAo8H37BwEs79aftEyzIM4wgVOj2bAWjTuPF
fhlSxKBWOKMIdBAaYeGIzlOCo5E7uBR7m097DuDH9uhinY3yESymVtwz8vLMKryTCyGPeAoJujuN
HFc6JjqzOmMaTpFgMVv2bYwWaIG2xKcJpzmWicajqE9sVIYuWBqDuBK/DL2nOs7vcqi2mM8LELfH
XI700eyf0JKfRUSvZQ28J/99F+Marxp9qbUKs9V3oxIh8rGaaEuunrl9f9VjqrAjApuH71Ay0f1/
JcoefiEOE9PQjPo1UdtO0pxhKf/nZniBI4CwR0W79pqWrf2pceOhaW7FaiohsKoiLlP4X+PjwPYb
kS6+waz4Fu3z1KDsJGiMDpYhL5wGxYRWiegOBXwGjSA4C/LVwExE6R5t1Oql8t/NIvWjZEJPVGpo
WwWCvr4CkmV6TpiTVNWyAvAte3lv6X7pLdUs7dyFwtd8jaNXHSY3hgPhcLkVue6NSfcXvbGUJznd
8vCyxoilcOkX+1sQHS2alazIEcEOd7E914V7noKML151hujB0ZkkSK4p0E+yYMhYhoUlKfHHBHpA
mxkcx0gqsthn5cJqGTXN0Ywm20FRJW/nu7cIKeWAWuT55FXu2kMyEu6oxxYfbA9Vtr2iYEMV81Y6
5Ha+gh3V0Lrxlmqztc6hPU6uulZvUcuMxz3UX+vPTC7GVxv0fc009IYU39EzGWRU9yt0vGlNYzeV
sGA+y3/DWHHL4270K2Ab6/oaj3Mn5H0dUQMKH1vtTNr+Z1k25QU1Slm17MuZrq6o+R4WCTOTtaUf
yO9uzGnc/QGY8XPWlorQqsJfOwEYzRj2b+9j05kgW4CaKwwDHOEmUL595RKOIiEH/mtYhp6JVdjz
eviWpskR/7Tw6//WLc0P6fdh64mCiWAKet1wfavbsBb6VCWoGqfqqhiVvGyMpQ3rdHeJXdwnleta
7tqcU0NZ4C2Tc4FXWgtnKohqNgyCcWRyg4UfLS2Ce1RzFDsMP0M4ajQZRtV6IK6HXBvjpdY3fUSB
CpKNgXzsE7GnB5FqfpjumSCowqDIQS1Tou9KjsYw4HKc8YmvE7JeS3UALAAeGo+P81sPuq2ryzMo
7z0er/R/2bjQ6HOC4DYfbKfvgUAj5pMhcqU+K/sQUoieodrKeTtlg/wkBJfwoiuZBoO9GZPYfpYV
x+DoMA3KXG5plHw0iULZVy+wypie+9zINhdBf775iTx83WNogxiLcrEd387n+TngdQ2DfUC6tDtm
AVO0v7vAXC9gub12RtPhT6uDYG5F5KCL6qOk7IrYhoD+a8fhuXOaxYsqbGjwDrGPZ+qc7PeXxsXU
oO8K0hJmMdjut3VFqtDHq2kA+1rPQ4KMyeW+9kk0rADKstTblT+Ek7pGKO/OWVJY6fXp53OlCeP/
de3hVH8AaIKh/1lU3FO3EbNxXbAzpLLnQGhdpsCt+QDnuYrhBsvrDg2jdwSx3is3N/sEnTk5+lhA
kudhZw802PZUnsDVcoO7LtoswSZTRLvCLO4qbUSBnCTkSuQb8eyh2rwcVNNQ+aXcmh7kgLUonGZi
2nLCBnH5YAg/J6Z3dm9weN37Nf9lXzqrgPXihAtEmbo3LanqEb068JtRg314kr7GL+oykw1J2fTm
HEE1ZoJe2l2EonPkPRldPS4gxZjUzRCO9lNB7iJPoc4vWpttgComqSBtLs2LjiZXcDnKT1B5VEFu
LG/cSna/nqdQovx2cAVvbUahx6+ePDyQyvP6SODiV08w3RujiLk+pOg3HGHvSSbtPxz394xZh63z
CUFD/MgxcRYNLX94fQ53hXmoE1uHsf/juHNw0swVvg9pKmECBXueEvHrnpbHYw37ENN+HgvUlmfW
ESO/qeEkeItfs9UtkyXLzGPDpbpAFK8vXghEo+Bas94fiwPbnron3gzRBcZiLAh1F1t2BTAk3QRQ
jfaR6maG67dXgT+g9pifYaUeuAGrOoqFc953ALlVTE7G0LJ05c1KnH43u7XgPa71Rc2JYvtFKHfB
vS8iyCJh0cIa+Ci0GoXHRGVTcytSlh9itXc20+3hRcK6WufzJ5HFcwsHplZ8oy9tXqyvV0GEiPVx
7hIBrwKhAcoAt6ASQ/iv/wbdMU691sQ3GkjF6NRmCS34F8nQNp9w0MGLkk51npCCxJkdN/gf2PXa
/jK66WiDuRZCbw/08aUes+GF2YVhdW6ae4hak/QRBS9d9OISiAtAPON6TK4Fa6YrVQdskQBsoxEw
peKG0DMZ/ARMGHz4cespdMFDvseML96ruVqI8hlDGEyc/eXikye/nl/Cf8aJeE5ITBOac2+fNPs1
DbHR9U+oWfjFNPIqytU8kSpGf9tsAwObLwmXaQC6vaS7rw4OBMntI+HFByVAe5AhFuaAVfmm/H9F
Ghr2/rp0p4WeADXmQf/ahP/40272T3ThiOcH18ztbguwrk99/IGtCS6MzPWMh0t5sOd4GCQ0znAn
KiUpeel5yYutaBTVbRLpNeDzcuZPwU857+0OuYwQ8PSCiYT1tNfzqDWdKJT7OKRcLLhNxadVvuQ7
bj+LNXOS4cA5r7kfIy0T/FYBW4ygV7hP4oi4AkHTmHm1bzq4jgfMQJU6nAL8L/0QJcQm8mcUtw/w
0jhqgt8SVn0Thl1NfUZkuCIgeAKUH2nRpO88mv3/RdgkeGZIfylpdqst3631h9tlCFvZ6RvJmyxn
cZtpPq180cgyznaqEC1hhxeCc5SouklBrO9qaFYFStjDnENs3L7pC4pJSjyOovHeu3pYKBmYlrd7
vKoqLxYlD57PI/M5vIF06GFQvR7ullh0SS8ZA7F1Yn7dcgKDLqojL871Vr5n8axxQ0lTLuPUIMyH
T88aEYcSMML+7z+wi4x4zB81VPjJOFfO7TUWATTDH/1lMSyzoJWW9GDRoNU9mfJuW27ohpESiN3p
ZueGA1kdJw16Dh5FG2JOnDjhYaInSioLUf2tc6I3+KTsP47wq6m2xQRlDz1NpnssWFEFLO9WD7D3
fAk6yN7IGex975iNP38hYj1EkPrjqyEIX9BNvU8dGusSujwgYZP33o8BnWwFkjL6/3/Citg4c4kH
bf5I4iKlCzm3LpMxm3pWuM0rqvFRSvcBvUY9NsnLaLONXwvgVGdyRzIidsZ5O703f4Ez3T/GtUoc
lmKex5mm1qzlVjmeXH2h+j0F/181zETTfGVaUyTCHALf6m8fnqB77oumqa2ID9y26YNM03L87u82
8ZlT08uSmFh93oyq2OEhBvlLQHRTZeF+/pzJUf1UB//LkMNNNgIb5t18bbqZKrsjor7uG1gOTgjj
VCeUyzmN82ruwIQobr3/3qJN+CT1dWVY3hle23DxhA0MHJoayUsK0kJ9NvrtkGl5mOa2gH1sSywB
/Q7jtVnCpukDkETtso67c4ttAhXIrtBGYvGP6enD1cIXJGJY0Bkf7R0Jmbv/U8CJvcRTaho70x2V
v3cFnf3Yhd2aABzzSHKiiV/VoJKYUFFhbw/DeRkJqXlxKmnpv6TFRCPdUqpmxzZF3Z/J645TUXGx
aZAa6UXJZ2NxS02/z9PPFmb9aCr5OR/tmtemsGqhWWx/jwyf2Qx5r+XLHLGjkTqXHHjjSr0u4eSH
cgWYRwHYjfR3LiIt0Fmk3d87ft3vRT8TfG6zMthGJd8ru4E47BvyMDfRnfI8qMpWlv5il/OK7Axb
GbKNitwXx8ogk5dJOtcK3a45Od770IkEn0SieVm63mjgxVsM5zptWSFbNgXt/h4a1OHN70Pt8wPW
9f4FLtrxSKPEQ1oaMlm0NiAXlWgvgyVejqfDY1LuJyOUjn9naKBNJ9fsODp7eobpeJDkNFk7XuD5
wz4I3dsmZf9Hbz4A7/9gLE6MYF2DuJz0x9GbwqVYAVviw0+q9FWO6Q42bUSXiXgPrq4vVU28EdSa
GJGjMhT8psXnUiHaOkRuZM127JOFE0WbQ+b+FlSn1CquwQi4dj1cGr0YMyGN+v+RnnbyR43deV2g
pDKf7Kz3ZzvtwiME0EcMkkOwYuLXw+bQNifItLAKD25OKhn1i+oqAWpHKxHAlLhj0qesUiqhBUjT
euCK918MbCNwnbjJHgvU8EKMHaS5exkq2UykRFRgB5cTjo+nSF17i2At+vJ33PnpG6EcdLnmNIyT
nrHJxbSYfmRO6E7NBBTg7r5EWHcNdB8HpdX/Xo8FrjpzKwvJJ1M1/uoAiMqsTgG5rsqUyhYU/Zoh
xwuQs6Kwp/blihUKRUlFw6NtpCwW7RIeBXu2gQ0GWk/A9LP/Pt+xtmQ1sSLVecP4n5ZvzOaKInT8
PpXcOAr4bjOFlHNNwKtOZtHGW7nsnVoQe7Sut7kTmh80x3tmbpZke5LB6o+FJLIQfXT9I5Z8oXGb
MuutCWWGahQfwuIk+rfwfw3wSo9+mtGNeXWtk8kM/85NCPXPKgo1p6W93U/YxgrVn2QlBHtijXKZ
f4///AAw/lwS/bQ0sfEjtGh5rih/lvPiogQSk45rj3HFDXJmgnGVec3Dflp+wIixVO0pDFZ6ZK6n
nNyFiaMsRnOnglEit7rAH3dQxni+dkdlthD5z8dQKu/6nCsi5uHOw5ajrdRGNeum1kageahGyQ63
mQRTgJbBDtS2T2PG75UONJYl14lmQT5aeTSzn9du/R+LlcGmHp6zmpm5uObI+RJHVaLgcNNa39ry
gbGZ7u1lTCjRy3TPfh1uoW5ObUqFPQOZVDpyw63VTZPgmwpTimPasu5fzKfqfsBqhJV9k+U81MZD
9MaUsT0MiJt1N5e2BpwoWeBCP4HxYmd71PsDtf5weRTUUUwZmnMwAJwMelB6a+7i8ufxLrQedPYM
mPWjS/sh8zmwGTIpFY8fIAVLEqDVCKzYVJa65UuQMEOg5CcDin1fN/1nBuTPcVdxWOoXOHbg/tYp
UDoKe10K/TtEG5lTwCg+4KHRq26qXuGLydgxH1cULlzEjq8olf4PG98cjONhH+wfLK8h4PB8DReu
xijZAYm9IXDm+GolzqrsCWQJ59eGZlxMJakeUVVMuzVGuJfYRkSetNEqeD27r/ntH3VOUfmFc6Pp
AmIvWLjC+KnyjIAO4GPT57SWIrdToON1kYozCgFXBCKjmXb2F3I7+DTtMN2uqugF02BhBGJCbDjd
WXlbm05vACIomw64LHmz2M/jZGga63wsk7mWrkBWKWsHfqkMkj1FSwBXfZ44HBCMs8EPOuRJab5o
N9209pqKvH9Z1ieQJxc7Gffq1OFUfqktAW8lmt50guVl+aSvT13Nmy95fCi8vR0aNL+rQfNIlAWG
0qX0KSqUl8XAGw6GMcbD9Rwekip4NlSoysl0u0zYJ/BcCZe/ScjsKmO0gnVks/NvU57ied0oIdHA
/AaOFXwnExC8e8RgT2C1qEUWLjvqQQzDyYqmlWwjBZKs/Ltg0XCMwEXdAhNsRyom3RIL5tsbhQm2
66utQwzj/gYzJW89ea6jww5CopLyP4k/p8uqGWxg1ZfJyS/iFqHWqlLdKZg9s4pDIOxdQj8D9Qvl
U//D1PiuMowXKma4+vvVuvKkAPyu8KiJRbQVUOppBAn6gOtmpYxQNq+MlgX32xo/UCdpOkDyV5KT
Pyr6DDHRQcG9VsJbDqgtFORF0Ze9vdijk9J3CuCA8Q8Cx2zYasFUyG9ZhiLyhWEa7bz8oeqbQq7G
ZVcLnW8CKAP980427XW32cCdtGSk3Y7CLNL+v970QqfUB3oX3U+Q+FTSAINtcdo05vrLGKseZapN
h7bSTBUhKFUq09ZCsvO8jgPND2arrL8OaYmbRdbfVM6GjA0u9KTBtBaCw5RQ35OU73cNiyUbuqK0
aFIMdUwNJ61v0FSB7/XF5eHtHSgTgmpBEn1ivfGQrULYPEEarikcyOpLKQIKkV6KV380m46Q6KnD
x6B6ItvvVUYhIqKtdWOy7xeqME41DzQQa03h74/cg/0/oCZi3zqb3v6Em75caePDON/zzYJf3/NS
MVANg2c2E++FCegk3gOyrpTBYA51dHdav67mLtAJ7qeyon1uHzyKFCpJoWUe74OmihJ/0mUuoSNO
SZNWnjUFjyoMwkDWHSA//z/yzbwIUP5ZLHVumtRyETtBdgKEtHRyIWcG5wIk/JG/lWxaBL1+sAB6
hZKKrRX87PxpJB5HyjpItVjHzUKuVey1hoOcUARQfoZsVgl4M0D9Yqoepi88z7TV49G3xR3Xzd6S
7I3OyNW9iVhwSF/4hDPlsg/GsFkXNXa2O1w+MuPZ02XDYECubewaix9m9Z9Q7bj3wJcqTvqxSbjW
DxhZ7nZY28LZUDMGsv1M9TwYZFINUGRpXD81LrhIs1ZhlALPYiWUhEvlbsuODkZo0Skq9SqJA2yf
L0H6J+zhQ/boDmjg/AlpPae+iwnOeR00bG8qU5Hz9fkaGu0rM74QJD+34cFhsr6JMBJMH3+5qIcd
bgosHitz/AyR93oTHIEQaT7XyFKFgnwLSzxLujCFpBFo7wBdZ3pZessIU5+Ahaq6O3WepH4Jt4CF
8+nouT9VzsP8BbfkCRReN0segqJ9+WgLvQVco0+lbzsGTt4eFudcPfgGQGnvuIhyBN/ufnKWuqbI
D/oPFou+ELVZ5XyiKc3hV7Xh/EkZ5tccEI6GUJymRfgV6R7YqtxxpWxBhL2XKQivD8pUkcwm9cF9
+v8DJtXFEQ2Ffja07BQUgJvJ34pwhxngVJYFVVLxYsqJti4bZB2P5ajQxeVUM5Z91eB/dJYQlCWj
yGS2V5DKL9/lgOwxBx6v6ixGcgai+r2Li4+kSTkxSZj8jKL/tMN1e46UqTYoRcbV9AYpD3tJhDd0
ibxC17x2HRGqvwxtHcmoXQ5vglOttMyh2G6WhvOqplKIbT9aEBCu7LLxanE0obmPzNKgZNPQU+Ir
C+IvMQ+Ooe0rps301wDSc4FtdXL9iPpzTj7XwsalZTxSzrp+7ASp0P9Oqk9uBDwulFxlSpReU1Pn
54nxVDb7FTG3OU1F5ZDAPd77kVc3sodUWtvsJ40zCOMqM3RygcHOy0sKE2H4pYHTII2ErQrX8NFX
v1Li37QtJ1Tj7HWExd+CUDFW2a3g3RLroNYzJgXs5RaZZFAP5IXNt8kedvzA28U+ViR7Ep+VvCRy
TlMIm6octm+aGBqkWQOA/PtzMsdQfgqq3Y89lR0XepBfSCYL/bRHkN0xIzbNB3oG+aNB0SE3m8y6
9hHZy8XjXbCaPgjDu4JQ9m/klE2mKSgRpn3/g1WjQ74B+0XnPALLYqI4ZQMA7Q5A7WGDdeBWAqr1
Ql7kZwPRbLfpD+y0YoTCBkv7eluHe5w24/oTJKsDtTT49XKkePMrmopUgl2u0SlmoemHbyWZIJzC
JaVUWtrSHZuHW02ZKPWQVDVEAV9rWGWekWrG97nc2x6PNcWvJiEju57CbmaGleLFkn8zV5zcfRJ9
KMttlRGAX8X+gAp2FQhIwn2mVYaA+wDVn1b5qKz/p+4u1+GO1hIUH2hggFfFTqQ6jR4NyBZdqHsB
MmEEBZHIneNbVAoHFG9wsl93Pw3PVibPid0w4L+KQeUD0WPcfgb1VwbPNI5KtERoy/iC2477w6uB
eMSlr+ujc8JCYWn3w9lrh+it4rZm9c/NWiQi60wqIcScCyKYRwbfbwsMSq0uhXjN0CoNJtCdpeGs
YxYtxOqPtah+MC6IaEdJEHXfbx2mxVWmZ2OpKZNysMadjcwpouraFkAaaNpXoS2vBSjJFkG6sFaU
rsbNZGz0tv0J67pMK3wnn2TLP8YzqyK/IapL5nJ9sHtr4fZVJplEKWhPd4aKBDcjXeMo7h4JPMH6
PC/rG/nCmGToz30HHpJaI0EHpDBMKK+7M1guxInbGPeC3ri/00vl9sRp+9zuEriwLqHzaz4yUnga
UL05wu/R2aSUOiLFCDJq9jQpnY5J2h3Kb8/uDJnwQ5YLfz0u2KewDKO7pu7jK8S520TuKrxjt93W
agWtsdrjXVT38UFsmeqI0xPnNiI1aFih2eF3rkCub1KBwlPE/+SqsWLLegD9cXVccvtbNSLi4zi/
e+ro8Rt+99lc3TWV+2xj4fKLRxYc0KAoJjMmwdeCRCmBQMwd1+rsaqaiuj0cpJFSXD/LVx+V918j
V4HEdy1Kt64fEE3UfKFjOFZhko/mhmOifgwJ+BRQe65ogvQbdpivNSxf+vF2kab6ZTigm7IcnZgQ
LHUmFPwDFqqaZ4sjP6MlYjlmgxKsMPkvKNfpvOHvN1epTycYwXbEHaVst6Hx1RWiY8DHfCRW7PT/
I6yGwMcIweVX1n626YGKcnEg8U7Jv6/WhjGR9FSMcMl8bYqkzEG5EpbpU0k5T6jH92NpILFKzcf8
CiLPDomPniqEInRLSQQOkKqN1yGghZ7EKL2EAhf1epUwaL7XzaEjQCszEwn+xuHCC2yfMSAtjifo
Xw1guAFlqr9eVVYE/8/OG76CpAMsDHsSKFe8LqDNIaqPMMSxpuH8up8uorNKv2gkEHwDK/10r057
xBFPwGE/fSNdYNQie5IBBKU/XFyN8MDdqS4m7GLQYyhg36qGav5ZFTXksz0+tXAzgposeuIAPRr3
6LM8Th1itgR34a0071nia+wSGQrP1wBBmwdUPAgPUMr9JFUu138KMWTAbIRWOroXTXqWlmMav0bh
uuBsp4HLLxtSbQPJrrGB9OQVmoWmgt+Suok7XqghCnJ4q+VlvKL+musxojV4G+djfqsRhSJoBefb
+gEAqiQ674oFk7GYhoNeb1D0B7wVPlPf9FbrY3xZ9ltQ4vvE6F7qeymA4enRGUAg1TsmadctgFmi
MdxT8Kal+53ikpvKnqCH5LVWLnwnEH1iYoxcHH2fZA26HfQ4p1X7WjnrEo/80aRRfNFImYhzFoer
ENao+g8LGRTVjArf7YJJjU7TJYWI8vEVbzRDc8ZR1XxAENApFlfhKCG844CIvRpYDfjAutDOGTS/
GCZ2yVMo8WvO4vAhJLy/PiXUNX3olqlLPrNMOrMNvWWwSHI2XxIkKV5lIM2KZxIAJipjnY3CiTzP
VtqKGXjIohSnR6ei6aiH73EdPXYBfrgLjphANWqciuavqfk2ULPOpVv0iWwfw20/+3Api1idRC87
lhY4bn4yF9gxHqOgDTV+7R4QbyAD2PHj41ZCKkiC8Z7pzqNMthjQB7c9fUoUjOYitCvqSw0ZbFLo
uuA13mJInUn97mWCNfChE3Tt7fB4QhVbEqrjPeSMWK8c59KrSE7kMCQVCXGp3A/x1+ZDtoNbtKJK
+tHljWO1cZkgr1tR7xEsR8CAV1Iee6n8+FSTOu7mXI253qlLUvllPXYpOgzNhKHXgI/Azc7SMcY6
TaZ2Fzb5iNMFGEdBYjnZ2oQsBAro7EYnpoGZmntU1MQlJIv/CAJgxR9Duj5ONqs7BGgt6I2ovmTM
ILAXfEqA2QS7AV0+tzyV7KsuKqGTNYTIl446ZQjYg4cITCJ7KoV/KGcPL/r2jbx10MUWDKiLc3cj
Na62ErdthuKMVT1mvwJ5qXuzjNxrMEqKqwm6pDPI5a0fQ+VjthFSU0kmvocPIfLR1Pkju+7kBZky
sZ0GQvhiGPMj9f9uzSSOs7FK+eJnHE1tIl21OOlbLbQDLAY8rXT5l/T31g+nN+4rfwwK2Wr7UJJM
+qYQDyH2mz0YaF7VvYDbgTxlIVo55WFZtZh7yqkG5NCvev6t+IFM/NrPP2lI7qSyjRqLA/ZJnOxh
WehtR+purFAyaEJ9T0fSX5u5nepKmvF/PFiS0M0WM0D5SXBNXx5CNsoKCtSUK4N87Y9m06Ph3Kqd
D3HF3fu3s4K9fl/VpM2nSogR9aB/wIfIbZWST/gbSNdn2QlgNhNYGq3epqbsNEOu+2KXzEqDeKqB
gYh5xClexCSkZQN5n8A2szTH73/J9/CQ5SusjURVSTEIFiHa9+twMqxPXfp2nnXBMUOTgYkVZE0+
1Zw9ooaujieJpRS5PP+8oINHy+GQ9XQIndrhZi3NHfQDVmRVin9Fekx/V4FWVt4DvWRrwg8WhY+Q
2BK0gdueGXd+mJIqPBAMGqqsv4y7rcA7A2q8X7a3vCe+xQsmWOXpB3m0yUPNoW1VUPoSZ1rLUp3z
IVWqdS9ujZQZFuLH+Iyz7GCXUJGIBAuv7R0G81vDNl2Kn2GTq9RiOXZA4C8xE5E0puKDjtzgkCA4
YW6Bk7PhAc4/c707Vs6Qy1NFw3Wtsk6au1Dlb9dqf4HUxMEuh9W5EuZcM/QcmqxDIUyp09NgTkcN
vsKtsD6zZcxWjXXRAYZ4/XQmEiCruCNj3CaZErLYhzM0XTICQCSscuopo6Of1DhR50MaM8WrCca1
K95KqpgAErm6APSXwH5FkevaD62cEYoxczrp/V6BZX14PgyzlgEErH1cOxvnGkwP/mwnxSwK14P6
XOuJSbwsU1APHlqo1RmYmKRjumLIeO1g5SCL+LJjT+hJKl4Bo8D1Lrc+F/lts6gew/FGeO8fhs7d
ktk5HVKPTme3dV59iJ6A0oTYi5XvbUm+lYd4J4d5At7JlvPCB9QreLE62v79UV3A0mq+ygZYs84q
+olxRDW2lMxCaw9s1IW0Hzz6FUzBwMS2gmBArAZqa5FV4dJ7yLvjqfDn+J9JVY5sBAMEkTrJfoiF
hU7/3EuxdANs+uKZMHPGlzKZkqX2GG2WmBfbzZDK0+lzJx6MBknw7Tiuu0kTyV3QYE8DYsEQgRgt
7HclucZwhEmxKqOAy0eLBEzSkfbcYDfMvBOk7HPKJMK0aEtiIy/I900c0UphykTXkKTaZXesIf3+
9nGjLr2F7X80BOJ/p7VWhEqzf3KTZy7Lf/f3MurrSEr1bA57ih9YuLgKoVoF8GsTHXyaLgwjxkIP
y4uKm9hr/37hjLf3KcS1fLhMKFDyUwzTJewExg1WSADMVMVxTuOXDAMOB7YUTR6bwnKCO35HQtxM
d7Sc2SmKEQkIvlbmrHAQvkiY12n1oFApEMk1oYqLL7va4JN+cvt+6prg9HyNlesoVRrtwi1egR0K
U1XM8pWExe8W7HpTJ2XgT3IN+hJNckBaJ3jSu94iAyaCQE8DnCEWI4JL9kdkjnD/v0Z7vcxhI8o8
a06KQjGNs+axzmCBAUWe3MYMJa/UnvPgBq6OhWQeOX/jCmEXl33pwsJ+sk+W7nP5lSzhrnzUnP3u
CBEh/SVfFcZOJYQvX6zhhMTGTSfa/Br/kum0DCxQmPWhM+CgZbgKAqYJ6RFacCVaTZZvM9Ip7H/6
oSrQLi8bwY4aSmejP3cDv8pB+cnwH9O5CFtMWB8rvUkQcjwJSHQ7N+NkqrrQkmDI6UT31aaMv9g0
MePZuWJ5QttmR1nRUmCjduvRCJBLbqNsDza/nmH358dqaQqpT9M5O5hXm0YfD7iymHrbdRypGHTY
e2J7bLmI2sE1Y1IC9JwVwrGSkE2wLAU4rkIDiovZDh2A0A41bzCh3gwvsIE5xsMxTVD9EVh5jUw6
7LJtZetSr+hGpLWfSqA/5GIvtHdqpEXW/DsccUqyTxSsOPyEdX2Nkno0T9XeW3YTqR7FJEZiY1EX
T3kzThHR8ZtzFOHM0C2rUX5UmS1bOJBi8XVAHud1XlpubocegDBJVI+zYbCBXGVTty6kLToCI/SG
RWXBpjBRsciecUjYIRSRBqsb8adCxfv6oV7cmRd4+6bruUSuH3Nb02bK4sXEIdfzwlX3kZJamD16
sk6XdfvlYvkHwuTvnqtKz4qjNnJgKt5FVCy2akeS26tySSD7SSBaHwyrt6PQ3P+lFqHlOAOH5qDf
5QCZ9BVFBKLLc5fXZkFEMNWfM1ffDIOLpGfjlMqQC2oFAdHj62tKAFGTSsznMUEhbBuTmCToIGDM
jQSkxW7rsFd/CFVjLA2ziAC5OAKxe36ezp7Hg+hnfBmmTSHW1PuRh57pSnH4QgczpSZw+jd3CQsQ
MLkvsrJDKaTjcBJr9wEn45NbdM6hIJ8pfWl+bcYAhqsVlwXC9bNyjk2xti4LUSU54c/H8qrd1xPW
JrrS8UhRhu/oxYrQ3/+fewRuoXGDqEcSXyUE7cH4eXhioAMQvoE1d+DCiB73gH+NrTV5y+HwDKua
jZeYGlj5rA/kLnJP8xtbc8LXz9Lb6ZGg/h77GxSqGc6h3bB/qH80HBlHgAEpB+DfE67iingzA7Bk
6CO3q/dOEXgRaZ+lXSINxBVKdGDwuRBk2sJJ1f8uSAx+rPQVbe+Drjhka5xcflED9e5MHE7jvGPK
vF7O8LGpYye0ICWzzkphz4fEWTgCShRueQbTvb3pzT07f9S4oJck4DvlZ5SlK5Ecdkef94HozdxR
xt4akmIDHmrhuARUyF9MMX77hX/u5ekanaxkYTx1xIBfngCCq2lGNBpz7nHUGw6aHDutPt675qH2
MmlClwr201MpcqYB/29heCrFbiOWd4NUJ2Fd7iZPQ8BlO6gSM+9cFyuLf34xv6D2KGApibMpSaXp
wb0R//bmBbjL4vqZaUQD3HBrIqOX57T/Vx3waEeYOyceyD+H/OpOAliqMl4ZngtxdjPZLcxYA1V5
aM/QxsgsB18YqN7I+CIL8kpD7zEWn4O8yIBj6DANaXFbC7EzAXEwSjSzFp3gY2AcRY0/c/eVLATN
r6cJNrkBvSJZSdRN4cUd8FsmWkvwRaClRRuK9PBP0AtPEpUkcFltu7gGMzO0W87JG91Dbm6d9+GC
SoDavRBPhmfCuXHZiopwSZGCpxaOSOXyPjrie6LCSkzjqbnrM6AY61vOnKAo+0SDGtZwBoN/aheD
TLva9/nDpj+rzm0Ym5EYUdEs1pQKVCKIKjsKwo5v0RtL+i14q4EBMRnlpSOg12vHIQA6PaFjBui8
lad7/LKuJ+hZudQP2IJsU/zDtSaB3jWQ20fg+rUK/bvbCohRKBLgpW9FmyKBOhXYYWgzszQEbmqL
rUtYC+haSjRjH1AWe4mTwZu8gXVbRW2ZIeKE2bqIXvTMlSBn9N8CS8f+leHRVhewb6tfGoHleOje
qIs4f78m9rMLJFUS2fMtWN9UlOyQ32eG4mKzq8OsVLzf/FJiVV4wyr849FRkUl/HrGCU2HNSPlih
kmcG5U3mxmYvx9TT26xhwtQn9bJQok95C4Qy9xSzJiKykpGnnUmjUKqsYoKt5M2K65Om5SXfoXnJ
pP+WCto2E0q1twPZtfrib/Ny6XM5LpOotGuCOAhaK5+GSAJACIwbe2x5inoBCdE8difagakMVZ9q
uk6HwTjL5SbQRsba2GiiAQCA/VhlnxwVjdm4z3hFm8Cq03HLiv7Vw9y7lGQG4X+7qfszWe9Z0+dx
01wlbu4yXd2otQZ+NQcE9bVWQlpUEj+N2aJS7kvpnvPa7o9rjOfxc+Y07Gjpc+GLWA4nAC3NyIxZ
mEvo9iuoulDliV6XoqVPzHD129DK3sxCNucqtUoaCzg3qOw31JJqAPx/N3UJIJxf0CVGbvWP0tjJ
SpBmdo2BfndTkCGxTSYNiulYR7Bb+yx7av+7BrpZCYcIA2bpgadoBx4jhrBwxucWvJxhkd97q+Ze
VQzeqg2BtmJ1tRLWqlmThzuPjXje09aeu26zUcd4ToG24ht0FrNE3Wi4YmQ+GlR2yPmJImciHhL7
ccvvw7HtDW1d+A81na1Pc3g5XxtZfNRIvix/13sKdWMCd3FckzyLrbxNEfsQVcsb3O16C7IlZzn6
Lez2wXJi1PJ6ubRyx6FYB92P2KIMl1IMFdw+e0/RCZsBjnEzjuTVrVQOCibMJR+Z6DTWqYopO46u
0xf30P/Q+VvmeBCB8Id6+MajY7Vbj6Jk1lXRB39AGvpYY/vGGIaI1oOINI1II2So0FobaSRCN0LF
UITxk0PsQg30xRru76acRMAC+YFnBiAuvowzBHbonHsI+VmuzRaYb/PD7sQcoryfo/jYpjTDDtRp
yME2fDVCdzT6OfjxgcpOJLSImL7xDlXbqe6WYfJ2xWyWBR+5+EeJ8ueLCLVjrawQxUxl2TzBXZ4a
Yx54Tnk54VbJVWL1Nq3adUnyyTP/F3UzXyW4i2g0a06E4ipvqPG91YH525pqXPjX7RC3bF6zqXdo
nHi+0+EOlP1KY6LOoiEnCzoPfjbGz268tF6UIB8dFqEj+YOdMZBrlnSf+Cvy5YiNYLQ7vi1/HbfP
Cua6iBRpI+6K80O4aAAgN57Uxpoo0r5DofbKxciigUsgXdP3KSZkeoIPjUEXW4n0rgyqwah8S9zn
pWVEbYQnBZ1Plpad/1kErPOKIFao4p6eOudS/RTGK1CDMYSBBqxJhlxq2mzB3gaOciedC8KRIqaY
aTgRe8aXRCp6W8pCXe+6C9hRYd5hQ0/pLJ6pl3B1aaGRKkDfVDxybmpr5i2tyoKwcShnC+PAgRho
4WgJBlP3svb3AZVRXKn9nmFCQk918j+SIUagykaxM27FaDR0YDZEBBkfm6IWGPvhJ93YSCzjKIhU
TS2dI7nP+xSUjAwVJaNk1fOY1MqqQOvXmnE615LvmSEoHuv+EwwgdNfott5fP2QCyqNApTiy6UR5
vZSg3q6Q4NY5ayVJvWrTWzr6DJi+dd9E7nsaA+aChXRCE1NaO+XnBlvfcZLo80uB3/DxyUfZrxS4
Y6KGKwzbMeu8XuBxRkMqNLp4IdMVPqDWB2t4QhI+mxeFxmuzRV2ZIbpsykL/1ye9MrkQaA398AGy
3j9piZ7gC9jH+uCzFL6wsOU/UklytlDPvjA0q7ItGAAoaEoyWF52F5vwk9AxA327maI0b85ip4JF
GCS8mUU4CeCuci/v1O3IjIo9Vmk5udlR89n2xHwdmzOHtQ7G1Skmgv1v6YpupnplzuONRyKuPBYy
Itkc6Q4KWN6DMKv8Ii796cT/2OExOTOlzO+UabYrOcyyW5ZuNg5zvBNlzrbaEF8TGkhzO4Uhs/Yw
nxp5EACb21MgVJt096A2XFC+OXpg1W8Tfmg5VAFpu/W74M6LqRVmkK9WUF6H1tEPN7eWwDIjO902
DtqD68oQlNajnvFWZngHf0Q/vKU/LJ3AnR80PrUqZR+M2qKnCgqb8eKccBMNwjx2vsAGKJT7GTGb
Yxnu35eHbpp4rJ2p6U6TgFUbOGiC3/3gmzVz0AtltJ4MR+Fb3W5c/3PoHGTjKg+aII95twRuDzy5
lg8ZQUI7u6Hy2/Vs+xUB22uS1rlFFl4jgUYE9XbKMl2M1Um9mA1EIK3W35uFzp2hiw14Sg1cYDJt
YeXwfIKrNknQG44jeupSp2vKrfawLNs9+xuRjnUP9WHEmyEmXmuBykl6drAKtrl1snYdTEEZYQEM
VsVOeU8Ad7IQDBIf9/P4r+OfLNywjovXvLJXy+jlqMHmwcn5HGUVm5Yp2IxzGM92rbIPAC1Uj/0+
V6srbZKgAYH3nMAqolZ+y0Y57C6PIMYHaJcY1Va85aPh7hKb28SMpixQqCD6ebAAxtWV8G7eMIt8
HynnCVzKm8jBT+gd8UKOU++G+zHsWMA+ypwBos8iXHGksw2EvITJHvRG3CNwHyJYYgnWYRCMb+3i
eCSmu2iICSq9CtuSXW2/HRXTXLfJKYj0lcIRunpyYZ0Ok4IUiWybsse/ii8RcVXPG5DDv+2L3aOH
PQOHg0B5A71XS7Xz3trcIb4mgGI3PkwWZIE/2tXPPZh/722y3dQH1QFubs3g717CgwesOl73Epkg
skgPDKXlem43snEDm9sf8EQrqN+VGFZT5hotG/tWA7gXeFYgXhIsimq0JCCUJszNaX4BYkt4s3d0
a3BH3FjWiq91sWqxCSJc0APfiKILfC34PxgBDBAsE+UY/Zm3B2VwNOVIne5jn8g8tbx1wXC4pPAh
DBUZgpCNp0rI2woD1pNvf5wzsBABENHNt3Csgt3qMDoAekkdDfkdkjOs6CJ0FFgAThsjVk1HZvfA
mYmu1cadFJAOwS1omRYGsxGo7oOSyoHhLO4KA/OhPzCYREbIYvXWAyALsiFgTclGUAJ/1aQMMpeK
KHUyMS9wi33jkC1e7ZfaKm6XsEsHMPJG7mVhFVi7EkqGAaAYQKLoOtoTw89PSwt616g/3fmaPUfk
yNd0Ov3UosfxSgfx9BOamRlfbzeL32VmO8y8AyBcZw9IDN+g9kybnCZaWISHUKiUYDM/j4s7xrqP
n0RbAtaJFrbbmorQeXe+Vpdvp8F0LcbrjZagEFAt45Qxyy/Jre1923AB+ria7RrG0mjIrFzk+1mi
c0HsunpmKqDNusj4+F4hVZpvX1u09qQ83f5y2qsBjygPv21P6b8yFn2X51d/ulCFyuVWTqxiKNom
Z9DXdff6ttjEw53RNCk65k0i2wP0W6iW6y60GEmbGTTmMSJtoL6XwTEHybQXjRxjfuZ3GKLcD03F
cdy7+yL5YC00AhqRqV5/6jiexMDYEg+vIe6+aeV446QVxYyqj9fmRu9fipcNwhFsZ17iLBpdTd52
V98b6tDLQdGcI8jw2Ln2uMMgx/2BKEqliEbYCN/irD9LQddFqniPr8Weznm8Ni1aeL+LeDbB7WlO
xHFxPz12CE/PL+0aMoWh6Ao/mqnHALyHfR5Cm8IV5dKA0ZhZS67pjacVCFWtZP8Lb3MIY1/lNGCG
m9yfyI8KrMytV3CslBOswf9JibiHbHYiY4Jb9REZet5KLcuCW24sSCUWMnGMNSP4SbH8UJFdpxdD
Pi9x0rmSBweUfqxvNxhO6hBMx7+9knRExOQvB2xW3UumfIlVJqRg25vRzCD7WTxfeAlWPmuLSF7Z
h7Ev9DB13zlDYUd5GbmRiiLtXgmN3PxHUG8sQXIAjyWSZepth1VXS1ca06CzmSVK3s1Qj+uof2Jg
K0zVB3cds6FjNhpxiHIw+3mWnqIXLwMrp9VYW60k27XhMtzMpNRQr3swMeaOZenfXcobrIlv1SYV
/z8zVtrD21rxFCtQWvQNZaMQmDlZKbCixi9ZQQVH8pLKCZHlVXLJRVkisL30sBTkfKLNmpxCqbG+
sBF5EGZzKWlSZsug119i3IvbYQbyYoyOWGGFmwrXUD+yBQ47PPPe1eBHA3inllHhpC3g2p/gjxBT
kBeD5ukZpWwL0ylsc3+WVbUxsbEDQBgYrk5J5kPMhICIDUnbWqUyj/8NG0DBbQVfIROE04MVftT9
NdznSPlmbVQzBqmjjS1XbhazZ1VzAAC65IjIm92ERtxD5l6P5QM8VG85gdH75vCpa8sEV5AOe5ux
Zqm7aR+Tu4Nb8zb3xfu2Oxl0/vLH7mC9xJvtT7MkfYKfm2KBUxiHHVWo3SI95lUgW91q3W4uycWD
1w/6jwLkJdA0D5/r16tFrd8hkEDClejlcRK9ivDM7Nr9GjEo1+0HB/g3aJDbavJ2zXyzNJ4ZTlWN
bBaajTGtQFJt7t+UDda8fFasLMxL+mKtpx0sb2Y8nvEIV/htXwKFSrZGPZ5iFDSWogvHw3GBEYEC
ivjVDtFUucMqLLH3JOcqLb0JoaI4cyJoDsc+pyUgQRmzw8HXYsIH8zH4eQ34Q6CkFsENj8gIPRYi
FJvCjAIJzIp2dXnFlNHNCFt9lFsG4PMyqZ+xjbTVr8R1i1vq5Q6MQdehCWZIJLh7ldW+JGxDNAum
AdYH0QApbo+JQ1hfLEV/ehaYCiqBIPZPpFfXhmp0hLPd0G3i8yDNVGrY9cGzbx+FcwURmSQqmQfW
72G7M7Yb/z+VFzA2okTx1aXW/0d3hJNnb8IjceGFDD88KU8RFyjmzM+tAY+ecVJaZJUZ5ayhoTru
pPDWGt1ZYrY4GS9Cdn6U64GqhS8ry0HCw11V0nBQP0jQTUN08RR40QQ1iMahArKPAPvJ+8x/kIa+
sNAErJ80xu9y+Y5UAe2jP4pZsCdJu+r1uLFlHenKiASQlm5BuDGQvILCVaZXG5xNADA24+qsxtnX
qhVboJ9XlbK0KoTS+0oBxD4eXyFG0H28GkgYEldZdvUWeH53/btpkQmjp0octY71jlSf+fpAIhMa
Ou+0UOdkEBTv5l47xpBZva9FJLAZ86fDsqymdpMBSTKkBeUrCov2nNv9KH/KIHiHdcKXAxt9HSvC
SICwDB5kEq/c+DHH/hLbCpbRZG1MZ+dz+xBgxrdCxKKdmn6BxTBjLYXzznmx5fQqc00Aqy8Lonsq
RIr7t79UATikRqD1nmft8e2se6pO+rz9D0d+//bfN52hoqulPAxgDnUr3F7ZVs2FkZmWCLURT9u2
PVdy/TAFjJFx7JtUr2N8x4Df2aC1NoO9isXHjejvIszqffYZRyi7dlorRbn038s2gEbqUwNImiue
sbWQf4r4lI4Cz/jai7JulkT/ecBdZn66PZtSDeZ68eJxq4Vzce0Z8ksTGMb8wbi0cM7G+ukcO1zg
UdvuCRF5MfluNRSRzyS+yEuKfawV74ELXZyrGN48TlQ7WtEbyBM6aVGVw0ssaEAvTbIkAeheRV+5
pA6lwY2UIV5l2HLhZycaoQsK6MgsCgQPIkh8c/nv9ZpzRTUv/PKRsA5+5QrN+An5OVBpytUIwigE
59NmEmRVJU2uykEPG2y5weW65uF1pXNnS0+t75zzKssFbwud/DZOMdGM91DvzFmhJWdAml0/oLD9
4CDtw2VDbrmLsc2/iMDx1w49XNaScHeEbm1V3Jq1E/w0UImVpH9Sf9hla+hHg21coQCB+kMC30uT
tm9+txjug4qLIqQCs6JS+L3eow/9QN8yl75Z1DMBtQl4e2+CjkxK6dREXA8/OtIw1A7h5n2SOrvv
TcE79ik0RUJyw8oPvBkZk6zEAHzn77oZT1l/LLaGsI0TCApoRffPM8JgARezcb2XDL0zX6HHsUQ7
TNqz1sS39MZuSXARc86mlfeD5kAUkB0OWgTBXBrviAaWPqFbgG5lR0o2bLjwl94QCyuw1bu1vYny
5e+ICGgXkninlbmPfju1LfrIP1kjh/1qvCSLiHf2SykhjZyHXojaM9CLLKpeyn3zWPTcuzY0Z/TU
1PJ5q+HguRcRnR3OJpgWMr6zhTFhgFZv7dpHOR4Kjl1VQ+GT27vMST/bpwh2qjpXhq8PCMl2/03x
ihOxll5q+p3ODW93YRvVao6wk7OTmiGwp3oo7lxCgIgbCrXoTKfF3v9kyDo34bQDNcIyHcRoxHeX
Pa2AZz3MP9v1dV97kE4XZ+U4+pSpKg+7d3+OZRnSbI+ccJCGp2JH8i4hfyqFsrnWn4BVW3WA4LDK
lJChRPNnHovmNzhNHSvHoNll7Lp9Pz/y3beea1KJcYHNxksJnTSMwr6ffNLPslGiMImUkJUMsARc
uOsSqNjcPunufxtRrhx3IugOWuch2LY/DH9tEBprbmzYG1SYUTFvIF4GvkKwyaU4eK/fWI/xFqih
U/zatV3i8KRZFbJTHpOPvdbUQjB10Sq5OYv6O+pVYXRdyZf4c+tjiM8M9BmyOBr8i1RMutZjnz6r
HTD5bT0wlzKWWhvbrBc/ejnbX9DlNyWt2WimLC1WqO1u4X3IHtNTUHsrH2w7WDGCZtwCmk/LkxQC
GciU7WNV3VG8IzWifjkbllaSrD8P2qjmRNdi+t1awFMqJlnxAygwcoGJyztJ5K6WlKFCaphijAz1
oWndx4LJE/l8SfvwmMNA+UunKOXkkulF1fsa6yKSt/0k+KjHsjb0wWXboJIEiQraOHZ/FrQ63jve
Zt531w/2TYFAv5pZjdG6rVagb5/dG/6ToMAXt7R2aARUzRwDPhctyRQg3Kp7lncmSWTxNqpUHdmB
BxI2d5nMte7DXVz/FAUyfMm0nTFAIY97/tOtFcRf5Fhkgq4R8dgXY1tnug2yijnY22nvuv1bhukw
3Zg/DD2/ZFH0zgylv8RqnBUjP9GJZ6LUKDwonzmcHp637F0BtdOrMSQbV5c7ujQ3G4wDmf8D4d96
wZCVBBogwxwplBuyogL5hhqwXtSN1hFC26pgegXfDhSq8MHOBbUyBRETl1w3mEyFIcujugwSaSM2
t3pVgFpa1RjK3YC05oqMhbRNF9//wsXb4Q0ugllUDRnh4eW2OFiclKetSMEOle7F9ivujdNt1nXC
GvIHope7o7bK7Mp25eNAY8rW6baQRAKf4pzJexEczt/tpfGi9fFt+Afzrnj3IHypSwE78sui9e9+
mvZqO0Rw+PJmBW98t/zkxH5NPp0NZVveH4RUw+c+RCqz5lmP0DfANLICekP+r/4XTM6nnlXBQXRR
qug24A5BMX08enCAJRH6/yKOSR/mKToUwz0pCrQcogaaSpAe5HLgUKo4m5RAdT+zgNPGInjsFrgz
2mN51vEl8WQQnto6T9DpR+kYzgRTBcsJAjgwd9pl0zjJbw7lWJpRU55wUbsoxgWn41PbmrXlVzJg
qt2JnFnWxpro1KlbP8DPdocsq3d+ONM1lsBCmMiK4pmAEOHCIA7TN0Pv082z1jbgswIRVuFQILCZ
EWaYWdTdvl4XhcE7vtPPXBKehPz3kb0vzhXM96JYKgB0Qc+o4DJdoJACkj4suLY3wTsa4Z67TH0x
ufuOZSjJVwZ2flVi4COatzHXMGiXo4EEBeCrq0SGRYgJZZcWDuUDD/0qTtlA9rv5upuaCtMNgF+I
7W6fLqOMNgVAzKS9wMtmMEnSRcxKnXQU0FFQ4bgCksbVNDXDFo+4Dnsm8sq9Ji8OeFJ/Da/IQfww
lpDVruIkQAsxFyUb0u7/W7DCdpjybZ28Dw6uVQiFcP3/NVGJXFmfdYoVMHTMZb6+4UcE4qTDz3Ci
bgCOXloUjsWv04YfXtBVXYf2vaGqyQU4KgDbCBJaxDqIH4o8oziH6X1lRSYP3yvkfiLVTBCNFCu9
xb4vi31syxSnKiyL5qMzZAKyCIvbtSUG7Fn++b05Pla4AFzMUUBXOKp0cyjjGq+KnrBILJgrbIWm
Vt11rak0FvDK9XnVwrHS3bgbxEmo7w0S7UBY7zzULzdb2RW8sD+UooG39RnBG1hoWf39L4QPy8KC
FvreLOptUP5xqH2Fypba4MUfhMGGjJi+s/0/D3senJckzs01PejY2ZeFMsU8Q35nTu4SQZ1Dfo6A
lJn4iK29QHwzq+vCJV9NrPkwFfv9Q4s+Eb7QnLT5WO0UYVAPPJpb261ueiJcJ15HmAfByiElsGIN
rq1kg+2OEF/G8pQuziV37EbnRZvBn5vwxBMAsbWPW3WRi1neaefDPw6U4X+lKKAsE5pW5g0Zjj0Z
TSjOI/aWGraJen+t215u799g13a5rTvDPO1pKko4nSPfB/G3RM83/rFb3EAUK8XBIbcs3oy78AjA
NvVCVBuV371Qulv7iQa0vvHMf5D/2LeG2MeKZTW7X1D8a5O9dOMccFA0fXacGZ5Zmj/SaSPtUw+l
aN3ta77Nj+AfYmkDCwYaBz1IXRR8Uw1JIQtlRsHsfamcNEK+BZLGZKkGGOgEjurEE/3SBlvVfYjO
C151wOCs+L6noCAIUQkPXIluZDrcSH1Q3aH0U3ttbqV7T9OCaRm/iFkPQj6F5LPh2sRep2ZtCH1e
fWF3pvC+oN/zI3rBZHfNu7bLZw519kkS2ELZx9pZVsk5SIatWdSKiDq4Geehv66zB5JedZN18URr
4TsNM/rONtov8a7Ffy9zEnRZOC6/EXj6lg5Z4LCssdywCwtn3P1pojWh/fla2NzqjxIqC627V/vu
jzwrTKveAfDKEytFkNzn5RVjmv7VaU4z5fRP/EftB9dG16+RGlgsy7nqdwSex77C+VhU0ClGBrah
cU5aWPsGMplgSMVtUlAPTd+RcVOv7GgSGVAnHTD9zgqVSFtuWZFbdN4o3g0f9vquJEu/iAKPO2Xo
QWkV9UIVutq3WkZIMtksgtYM0nKutVQEgaA52bbEEsXOkx8DuLqQvWLITc4QB+kG8w7LJJa/rr4U
cdRxiwe1JbGGQBU37NLk8W42TwD+2K/5UcX6JPD8OCr6lzfBv18qujUcmKqxFZSMXrYEFCLYsVMt
F1QRDjONY7JvP4d5xVLNwJWIQ0Id1wTwL3ONfLmKq9gNaRIiNI79415x9MUMDeBLdOA8lVfZ0rN4
TPHlBIF7fmgTcasmAoGqG6NJT4VMpP8GWTz+aucoFOfdNQp+Th3Z9BYO1ZcRrlSO+yFPqs9iDtBj
O6vDDc8kEG5OKATCHmdhqKs/BkiJ7BbQ2026P+V8HZcmf8+fzXHHl7k8WbzlIjvlg3RlWFohWqBq
D3HHLpKslQ963zeD3S0fzYkGa9rOS8ujvWN9N/XPDPRMVNRnzJR6Cg27ALAVE6c+mCntdgog5qju
z/0C6AHF0m5ozNNp/vBin+j4bbFrdpda2AV2e4PnLsDeuGJG5jedmWFwaq91mrNmjQczSNPwIOL7
KaPjqwBljBp6Yzw4PX3pKUv32z+UyjCasK6ELo7GsiPwsVRLW121g+K0uSVdd/pEqSTted790nrB
guO1Wm2dSheKpeuJNKCqm6py175bf4AVRjAncdTslcRELZySs0T+ttHEaSHWsJA2a7x2WwPivDuN
/PpDJuMJbup2Or0NrM7F8qzqPBlhqXjjq99BrRxk9wYdVZtUXFmLPwApciUl/TTHMpaDr27Z0e73
Ra0csFCeLoN7+hp8T6wFiT4AE5GjzAoAkT+VJMR0gBAVaXOUqXSdZlCs1yehJuj4XIyPcDCLMJXU
mcba3uz+j66JZPdR9rN7BUMv0RH7Gm7c/Xo01o3LmPaNCsLreEcbl347LDuWzQ7e4wMgP5uC2TrW
Lq4K8XhkDcBpEFJ/40J/YvXjYidl+cGgUxwe/oEELdX4eDrbVBc85sJFZkt5QODdJUnEHeUaVJo/
7FFCYADE46BVnrMeafr/OaAK/XN7GrQuuxfOfnenLo4Zdp1Cjr/mTVGiwV+xcEWpfnk+Q0sEQAZq
curk2Bf6tR5TQ7KDSVZ233w64RivKCDU5BAy7OzGwOrBuSm2a7G+eX36x8DxsQ+IvAx2e5ckNzlH
Yblr7JNA4nhVVCje+hJRhtBV4nz9RWywGAUdJnV57Oi1FyovzZzYBPWV4+3cgYqgoFLmPRuseyR6
OIN29BD42coRjl+poDK2EmwHVsoo23QIQq2B6xKDEQmccV6F4AWm9kmffZ/R2b/asUoGN4TBLcRO
G0vjIf45D+thE0iO3nKu08NaII2sUeXZ67smzhZb64Je50MknTH/7HArp4lOfthW0yPe6pcjlNtV
yzBJv9ExE+69R5ZWVhns5mtWbTXztLxC53Mr+taVLFmr6Syy7R1sDMI4T2yq1r5DhvD60agEMsDN
ZqqvOooOvF4Nx9Fpd1lOSNOmYT3jMXEGiCc09/wSwZBFfRCR7fZBdp+0qnr72gyi/hS7kasSPGs/
sOtAPY8Fw4tWWw0OXbA64vMlWKZ5HMh9Ezs8O88isKI5Qdz0dg2z74iNckhhaUZXHFuA+bewA/rA
UmuPZucSsq6wk4/g3OWnnZ8/sviX30X6vtmMsurZDGjzZl1dJaQIdjObbJvEDS7mi5cJQPoCg+dt
55UNsPzqI9182OU76jrQHNd01YcH1UuvUlmOmbf+wbOcsAe/2tGuOF/mck2gFO/hm17Sr5PkKlzc
hvv9udQUPn3xzJtyzDlw+ebqNgmaxDX222qgKsQ5joI0bLOyHNWMTwD6sHfEENF6I5UxxWfM7RRz
hQMfRWfoaVZMKLfHYXbGXREVgscY/tUON8xYEl6GDz3ufrm5RqT96ZZRKIC/X7t2u4q7jpY+lF9g
u+CVoPiliRdBLOpJOMCdggoP+wN3KKiuvTMmaDIDoZaLVZOa1O2+V0Nd5pADmB1b2UtIuHGUuZKO
nf1lHdb7MCu6n6tal7uFPyvy7k79lH4B039Q5VPalsKcKMXWJ8guvRSGtxyn12x73cC5A8IPaygI
CM3iFeBi3qFauywNtLf2kpWrZgWiFrirnzzqtFyVYf/7Vr4cMPnZ8AGPFSbNmccTklgy5N7TnQlv
BMNAA9XH5XaOMcsb+SGzEXwyvKJQmmHu8b0bHfsYH2r2+nhGcfoCRNyMiscqrrjqHLLhKRe1gqcw
llLKeUirWpWMQnDI2oNbqovpflhgac77bz2nFR3i5G/RAPDW/3vVvY88J44QA2RIahAhvVG0W0tM
6QOoDzTjRLaE6NGM+dZ6g5XXpDe2FPGWrllz79jwGMeyCxTSMpw3NDOJrzhisXIEMJr6xivpi6fK
0uFPA3bb9svX7c5YjIp2OoMhC67VxcSsgpRdPxfL93xytc3dPbcqLAUTQv+0fTtObUATtVEyinVt
xN61+uNE6MlYnj06nCYme9q3915gsqOc+xw99kVg98k0wRjLb5JxJ4lFlSTVERxMF0n4KuTuWIeb
sdIHTrfnrbmrcHT4pEanbtavqZnboP5kDFDUZ7tAsN3lktrEkO7mKbC9o+f1dL+BC61N350GDyjO
cTrbsbuQfbjV/NvFWmXyFkc1P6DCj7Ei88PqL0VrS4oH0iv/L2BxUvnzXJHjhOBSHzLbqmpla9yp
tJTnDHY9astvzdqiE4uen8lu83WCf4UTr8VL2NpzaVzze+cW/KFDYSPuVz0I82TvW2elcu6uTV1q
KoRPp7WBhcSAfdREbrB8JkfEJcwKPEAM+PwldWkZbS+UUDLDAO/wx6cYlNsAhVHHUqu5JSkLRR/G
XCZW+mxHvxVT5WR5iGy6GI+Q3v1se2UbQG2s6UVLk8nKeWCmYkryJuRLHSfcSaAs6Gv4EtFJ80dV
soaslxxf/BCrbYFWClwMNfvgM9MU7MlCKsJjDNc+6mJ/d0MLGwmok4/xYg4CwzoRkmD0B6TL0I2D
P5duKg59sIVAmCTmbmDHckwIqXdDKc7O4UFTgYfOpfl/gAekYoq5JK7UQdBX5Ug+vVyIwI+Z0dbb
IXXNxiIv+iKeNXsQ+usgOSao3dwSfAKcB9IPd1UJU8wQMVgrAEaVasx8knnu2ZrdSuBZWFGZAACU
j+Nw8cOUQ8nU4fZ0IAgGRgq2clZn1SWeKFqrwzy56ithv6SeW7bpSBRTZIPiBnUpWVY/j1jtgXqZ
TNz33RZK7RRZdKBzZrRmKZu/cDFlBdXHSR7V9oE8J061vzpuIEh5vnfQxPhx6LoZXKbZRGTQFNZj
kihBMPDd5uvcrn+Bc67iG8wYiYIcMKVoulVzz1xUQCguRh7IPPEFhAtLOcsL4ZPVbg+80Q/S2RTX
ydNuwu7HZoMDCH09isGSFtwYEygvsTz56SHAz3kIesz1ghKZknrPpYIJbJV9oH4kLdcxQ7qUGD18
THZdxiPytvmey8oCAOy6iVqel4kuCItqD8TeXkjMBA6WbF2eZQ0ju3ridl85wUXSfLyOPyv/iKQ5
RXjgeHv8atxf1gF9wi24MuvgZYmV+6selJS+W0gH6OTFGnCW86P3hp3+Wypo1IBZuG2hBw1EMjO0
1T+dlRmEDuASPF2qqq7GkQmGWxJB+xnQ3Nidq9b/W6JSBM++jL/vn2YCuaNOZ1ItDm7UEo5+EL6Z
xQrTyTpqgr1QUx5SeuFyaRGHaW00OvzOxo1PLCjzw5yBHZ94p4/RcO2rtrjBFd+C0eruc+O5BWMK
C8JlNR1d+EVokW94W/Yz+Z/2bcNRd416MCLzJ5MXvvRJLWZOFdVU9wY0RmMAgDpbTr/W1xBrj4Ew
VG4pLVugAhOExiDz5GgaBSJkdutcP/Tb3egqYFAVOdFxylP1ivGe5y81kXHtuAlUKkZdzUW4B7dP
NHBNuade9xJUgTxREPX5dlzT5dWy3PYbH1NvZeMGxcjTuN1g0Jf2rQKBH/ODsLz8uexWjueoXOUL
Ax5QRiK5I9GRNnZIz3Tsm7ktfme1o86cvZJy1Pv8jJ7CHZX4dRtbx2cdhxRs4gM2nMrIIqVgL7dL
ck1GfOVKPTwKMdKibJFWb5WTTqFEJ5rgZWO7a1QtnI/Ry279d3BaxvIsn9as0W7WTOOmpJHp5FZq
SlNOUmKcFPn1OVUaN8Fsythz9wbA7fbKloehPuiU+x1cEnSVLrsLiSTNN4C1DZunw5N7nOBhW0oZ
fTCO57uBa9pqq285slu9MmHQva0SzWgo+c90skwmLfr3NqEZLPBdQ6P6DnocsGoYs0Q7rESesDig
rQjpkTLxCXdahKZ9th6De5U3X/U1CpSMNFQPTguSCnLj0CKoLt6+IUnpeiQ6+MoMh7Wkz8uh1b/k
0uj6ODKGXlbXy14BC34J5FmEFFWgeoxDIh7+HVCZW2Z2lRfvrh4yrZ0M7WnjIsN0sUa3yclvbCI7
3Rt2Txhbzk5+ZLRbd2Wnv0eBSolCaEW+VOxEQBjf5HgIkZkUx7r9TtOtOeoDA7QJveVQ1H505uja
7Wqy057tAqPEcRXNZttFD/7MbIzXD7HQpYlVRXgOUwkTKPFWyJgcOOAjZAZRw8nsxnVyEgYk0Bzq
bVvpY1eyB3jylhEJnZB4w8QJxh8xB8OEZFF4TY+lX2XRH6lEkjz6WZNvLTfhiVTY+1zKxNmB+OTl
2GEU9xKMxQAfMBk73YK05/gzkhC4FGZTLlgBmdBj6fP1vC+UTAVsUlYSczYY7GLBUU5qAtlaegV3
Pp9Ys1+JpGxcbZgOZBwLMWK+fn6w95NXzhcZ+YGGLJzHZWhwJEY0CueolkqSlfcfRvldwOkOpUg5
S4eQQ8Mdzhbfo71a08QK9M8kNpRa5B/Ulg2GwcRt4g9W0NBwjyGWm4lXwn1/90lnZQcb0RTp8hvj
Z37FEh7PtYPRtpuwV6+eHeVA8FIDObJVnfamJ5HP532vaGNHsJiNIGw/fcsbqfyI7PtfURVlfYZJ
P5TZqyk14f6r3WMz8CCaN3Jvf/4k8W85XSS+eiM3WPDSHBudLYm45d0Ma0Okhcdc6J4/2FJgVeg9
LdBjn3Ho+hZXouU0ViQJoIy+1M3OfNdXzygP5N/pUjC9u9KG8pd//xHVxY2zM+FAl3Y/SpeB94IR
lKve+9+qZzHZWT0LzIeFMIDBKv54JHo9h95Nh501aGuelgQZnrsg1Oi5z2zv0wf1CYoBSyg5Lilq
MAEoRSCN1iUwDVx50j8KjabKjjNmncRyK25oKy885mYOciYGmCCPozd3FPMiDKUd7fdWifio4h80
hDWiFgQJEWfWiWHJ9+2AyMETtIZhIkyDETqACWIqQVwzIkhLdaTtBNGfOPplJy4wiVP1wbfODTK+
E9sYBehxCN2FP1ytxT5t4cA9nJt7aH4TMluPKQHhikQWcDly4rTJSjhLHsRtVt5cRI2VFA8eUvkA
ysTZi5OvLpBeiDg8+2wtNOaOFsiRdPJ5lV9ZzHgDafnCoDFAexmLJSp7cm/WWuQN3bVMe4XA/89f
797B6GvWv196rqfW+ZYNkUhhSmBC7F4j+3z8e0l/HautxNnLgyZ4GUyxHodSjSxdzxSqxSgljxSv
Orlug0NXiOu+3xL3c/1du4rtxyfRLAqxCCU959jcj3rq5DAA/VaGMLEQT+U+O+oOfTcgo5EUsJWp
N7x7OFR4cmoQgwZn6S4OWr7FEG5R0q//1wOn7uFZQ+by0+vsnWnKQRZSer4E60c3gy1J1K0ONmeF
57XyF1uIw7a+TqMrvFQYEHml29AAvYoKp/RsZSaOeW3ZjCWpPep6XKZo8Zd4aShlv11uhCsa75ah
yYAInn78pjcplCZ3rYqqdnDgkMs++sdrfQeyIOWUgsQrev+L/KDeBuohkGLENCmoj4dKOJ61BynD
n8FhUKR9yG6djmFXGDnuf8Zeilfmy8GVxLaJd6RP47oA/YzNaL9oqCQHbK7Sx2z6RoPwdozuNOPn
JJUGUig145I63wZaJof+mKCSVqpBqXgOkHjEb6InJhMnqBhMGnBvPPQlmwiEY3RNr/ZLBUE61M7z
hn/gV+GUk9o+Ck8h7ztnuuBddlPp+crATCHklJVXqVH88i/Nj9QhwWLDdFl1VcnP0AFLMC1MISCH
MehNQQoKkVomWVawXKZAf/Kl0tFPm33ABvSJRo3T33fbqOFEo+3pTDgpWJ0hBPANVD+25zpmuMgD
SyLqc4SuT4zVc74hlDRE6f2A/OKBPfRrusbZRjD4K2TJCPtccnqgJZtFg+fCiyv7FbRBD36Qzyev
IYrjrIyMojS73ttt3pt3yHsKaLD53hiZQNfntnf6Y+ismyeSrDfWbg8V2I1WbRCy4jag2mc+O+zC
iuirwAxptdvco/oDbXYaLsqo5n3wrTfvv0LlF32/PRRn1hs6SeyGtFxEs8+Ky4YHnX/gTfMIFmkF
Dfvhqn2kZaU3Z8GhlaFDbPRBnWXRaKj21PoQzugCkhFGw74/dEY+4I57CynXN9Fhu7/CbcwO5qA5
/18ZlgJ1yCpGcbEos5boP5EkQaZ+soVCHJNpBi2jv1JNs3DwkxCKtV2ACWxxMTIWsVea2ekXHV0P
R2Tymi+bael9gaqXpgFFXGKipYOozuyva6v3iEa2in/UjI873+X+eyMe1ev9EL9ktq0hT21NEPhg
jXJ4KrLJPO6sBUux9kZKX1K4cK7J0Xm0K24jGOWDQckkTAXPuvxcq8bjvAsXzu6UdYsu7hZIw+Ai
wGeF8/y+u/eZsutJDmMpNf3nDe/vhe261BByo/P783u4rBeJwXC1yCRlqnpiwC+eSzJVXjnN3nku
JPriQF/X+ldVPMf/6N64iUZfZhis+0MRl7lX2xkUlCfY6tcZ9p64ZLdLgar+zvcwV3HtROERx1wG
2yRono8f+gaWN+FnocayDSlYSq1S9+1kPGp07o6SWtt4eLZm0U9OCBCn8VT7mtyugQtR3oxGjcNM
WW7wmQpXpyZLByCkLTwu8EYggeiaS1pWV6JyOwxrNzOKzxxTaALGK5Yt1XxpH2VoC5j2HX8G83x0
tN6T5m/Hx5SJw3fvxSy45dH8Yp30SlRfxedLlx3j3PAZVzU0q6amMV6ncNjzytSdlZoDjHnJlAcH
De0Zh1yFWhfRueDp2i7PYz0WSqv+2SpoEslT6qNx4TYGdvU5Y7J7C8ZArCHjT/EqxggcGgpWyQvq
JZqZao4bPwt1tDTyAeDX71bh6HxWBj0DMFkM7wKyKp1AQkD51hvCfeRK0kbh+GId4sHzu+i0AC8B
AFPl74EEELKwON8ld1q4FpJXoK2PXo2eHORQ8/6mIS3CWfpPSyU78RTDhPbYXlSVg5Z7bU7SP2zx
gAWJ9M0rT7QfYG6U/4K229POGUq/WsfRKDZRRp5ec/DwrGTfCoGWDflpTmutKMLPlegPDT0lm5C1
21VdWe727uIx40kjQbkk5JYYig9lKt4lkgRWytp9Wp3KKlP0zqmYsJMh/DUASmPAi3b/4hGXd/YN
EQRHF4ey++ji1dxRkcgSAmNIeRlXHfQdG8I1+x5HposSsZjG4TnLE5Val4bAZASkvylRoqXZ18Er
CCyd4/XEAge8o/ZJr26dXpICJlE1JN+wovkAjMU+wf7uMu2aduxtX/8I+oluB5/RyFe6dRn/iylL
w6AMNTVqCrRzaMOPOaaiPJ8QAsEchdVlfe6DEdPi4M7OnZIP9ciqDYUWfsBh+bdpSlxaAbB3mwiW
DzVAsn1aknZUM95z12gnl+nqbPEGVDuWxhbPeHTb2yh8/ZZEjHvfdJSxeevm93qCslw/vLRjuPCL
XlAIR07a6tgkZ+gQV3OIEHayyN70pBe2to8L2wpZTlf/1dNDGYOcYSGzW82cKv09aiSRm28yDhnj
wgYCUkim/PPMuhQFboMOqGJjn5Ekgrjv7JIZocwSiI5Y73/c/4kVYITGGgIPgJqQSAor2jrjjKTm
8s75q7agYAMdqpbjE0nKb+O3haDJGmMsxUCyTY8bSFp4qtOGCMko/ujBjcABfZAMrXOOvshUXwv4
WvnhG+BPQxb9tM6pMG1xsdtpIkGG5hTkgAJwUy+3Bru0vrRbfO9EHII2TkLU6Ck1EXCgWVqt5/0c
pwSSS4cD52678y9MdMXwhugpvwMg+yyoj16bQFE1bMWz4ZQ9B63h+jdVoKm1ACdLjm98e+8WxBEW
GJfHWRRxw5PZITh2Lc8158BfTyXrpHng2PWBRhXCToNrPzjpaVeoqh+Eh51/iUQ+i9bwRVmihVgy
Gd8eGuHAIGoq0UTRoViTu7s8nrLbpAfaEH6KWrqlJIhGZ1fuC/3D5s/DcmY04e7o4SfQFMo3T4n8
LSOKAyCfuZ5z7QLSBdwiCXopCT6QeBVpF8fKve9aOEauRxi479eMTv+YW2E7P5q7j4GuQTzk+7lr
i86nAt7QqrWgoex6IVxYtf96YfAYMXHjFlvp7mMNdyYgLoCCr+MRXtGrjrlIvy+vPEu4OZ2JfGH6
5SLqez5TllXOaUKtEx3eG0vwxoRA4QF2LNb9bOyc3oTzY32jvrh1g1bm4HfdMrODx32UlMoOzu4O
UlZY1Wvz0fbKOdOOWKqwt80BYZyPnmZrRNSkdzc/M030ARZn/OcLNVSP8Ghf7OAvH29mWPxz+l8H
DvPPv7pzhI+Cxk9qaKDV2nw0UHF907d6uv6O2G7+7Jzv4ls1pW1lLNc0A4Uo7FMF9QV7EhTz95aB
3XYQTawMqWuIvClADpm/s/JZ8n2qRiv3Ubl15bDs/+lq2v/c+2h0ji/CxN0qhPE7DwF/TwtnbTc3
iVJNU4i9mmzf9SiAbdnWyD6D0mdnk5umU2l+KrX+6aR3NrTdPZbb7faZlMWmN7+bv/xuveNr1vHk
2fG/wquv4JXOWJ3xeMmhluNWO0eyk0wHKsTSVdAaXynIu6MLq0tUocpn4ehCbYJw2Wl0chdgQdks
xg0Wp0oLoXYU7ZpovjnyeOYztgSNc9PEOk4PIrxPz90omJVsHcOnbPV5q9VZT1DNDmyjW3v0c5vR
7OmDczG1e2eCIBp5SL2/+2IcSPFPLjhe7Ail5BNW/YA/YAdE07bnBiPDGFilaDghXaP5DRzVCxk+
OyTukt2+2hCWtVPZ0xP9afFNDWdpXaphhiDoCfaQlxPQCfWNgMjvsNpftVTSlBa0TTmh8A6suxQT
uz90B0u05YYCOdBPzSc5eFPTkDplNn7LwL34PMKhsWrJzKUWnZK7HCSKmW1+0kC2NTHE++8snON3
Ux8KlkagiUYDN05s1dwfVRQBvWlOuVhM20S+Md59u78bjihLQdSTWbmhhtSeAGSzL7FcGvmhO8u0
heDiJ4jm2yT/jHsIM/BJ8TB2QAEWRhG6SXZtGaDoOr4z+bxi9L+MNaV1vyk0mi5O4eCUKvQ3uv7h
f/5/vmJmad3F6/WIvsZyTOMgbxCB5l7vvBcGUwNOobi9k7MVie4YdEBsNT4E+x1//GzhB3UoVvbu
eSQ0Yraryr3iQahaGY0L1VaEzQZ+F/m0JoDNP50fkkvevgW0tyH+e45rNJmG89lDHr/fgre/y2ry
Po+iqG7q0tHj+a0bCS3vyGlMBcM+l+0DH7B5REw+ZFJlx+tBVO8upvkKGwrWB1ToVf9b/uGH10R7
Zk+ohsnkdgYRE0uTkEB4HnFcikXDjYlAI0/YJoPSE9AhDNBkCUu17QJ2jFTWXJu77gLNnzyMoNIx
aypzIJpd/6qZvtjX09X6rqhNWeaP+mv7aLp5T25K4ynKUq1QW+MzDwCikdbB/1B7hmhqLdqtse1b
7QcWfvwpnR1CkqRFzn2g7V0D343i+vX9OHJ8pkPHLL9x5SRyz/ngWZ+ftD8aP5c4F2vUmllCumR3
+tDQM98VsW/+VcS1NqOcuJUHl34EDLLQe59qpupHXqg5+lT7x5Ul6k7bPLdvYF8haIGoaLIHTOTx
JE0Vw1Lmw4yGLyOWBf4Q0iQ4fyDfBRqra5qeYZtNuNsvvjCq1gB0UCGNFMdTCpnEqyWlCMnAU0Hy
Ez6JDRrvvlolAzx6uRqkXAHm/9tsvuKbqsW5dVTicVWD+QTFFmiwQCkjcbJiPwCrsndQ9GpRmgP6
OHY1XE/CUWs4a5HQsMVK9OvbFrCSzisduk8mPAEneZIB7CSjal59Y8YVjnQdW0Gac+aokS1F5ppc
JHZdCmH9cWTaxncY+gFCP6uMY+Hxj8gxl9KMKk9wznBEQ1Rxu6YIxMTmY3WdDy4irg1clCMDU20A
OfvwT5dvLk0kiuPYKGHV2NPXWW81z9eIgXSFMdGU/2IekMkjpQNTFQklqcQWblDU95g0azcIQ7pW
VlELjvEAm/tvBaYkPHbT/ZnZdZNrNc3j3YGOY37G0CzToV3/qJxkARCbIWjPeIDOdgvWj87/T6RA
bIwA63XYdr0Dd/S4vqOg7FRz/LTvQMDbtqpNEnQl36EahE3PgOB+cgqK5dKbCzWB6Z2sU0uIoJKA
uQqNfPtG2yk4BJ8yRXKXVeGjGtb/b/NLugXnLRHUgg2HnB7cHEaotyjk0vYjFCrEiZpXoTSbntQr
yKDZdwV/1TxEd6n2rTyXH7meJHxZDy06PWDEpMGcZB2fJ/Ay9OPEyotg3DU0hEMjgjAu3TmLBH0t
u48ZmtEV1K9xe7aFIdCZe00OlO45wHYz6GiYajQRjMO9q7B6kB10LJ0ck/80Q/MvnQ+UjC3Vh+fc
uJXCptowcgpDOHD/ckbP3O35Wd+E5vTRLtpwTAwcr5aaGtOedIgh/tfwJ31uXc9OByioHY13rgux
mwVHEj0xuUlLYyaH7dEc/CaNNbN7lBykc7MS1ROuTGtaOkfyZOEJ1XY1lSaKHc3ZICelHuISi2sJ
UcAt2i+p1k+hJJ31UzLTkQ8i1vbr1109wCdWLfM/c/EGlNgCpWehAlO7WOEJAh3Da8YpcugMevqZ
bYJrSlaMO9Ayp/r9Fue1LE0Fz1lsAKlB9cpUwSwY/sn6/2hb1VUD9k1erFFauULNHDFThyIYkwkX
NsGTVEDHuG4XtmDqMzGdRqTwqb0/OM0l1LrWRMwHRvaOEhq+7aiX4UT44RvoIsRqp9p0JREr6oba
YZ4NlwntVhb105HQ8NCMFmXptIylvykxN1ufhc9/EP3DAoTP5mT7EOvxinqr0yv3Mb6BRP076XXK
XkQ9uqOJArfrjpiy/KBa9fSzh92bQ54RhOFRhTTGXal+qTyElY/1Zp8wjO++8bJzM5dzlqpIalOH
IzCHvl4MFoUgVbe0K1QUZ8zeN9NY4VwxnWBtxiEZR8p2P0eE+FdSWsLLpJtIsVz0iDQ262IQmgQt
VxIARfqIz1cnG+yEa5OhiCwZWTgxX0lSp4zYVfmzqMb7M3O++DvMdDKxZx0C3r4OPQp//pbiP57v
i+ln5Rrdi+G/fOMxOxoKnpBVvtGaXyeQSEpbxuVQwezuYZjgWMmsSpCbPpAY8DoWszupDzeUDYp8
/yqol5iQ2s4Z5WGI/JSjKmDwItvBrTV71eq4XE9+pWG6Z41Y/ucSgfvY/ELVV1UxsB0r5velwfg9
HrYh1vNrizFfk92pBGhbhqUYLMzXb9oHORHNWJJp1MomO2ruSbLMEok2eTTCWHdQUHE3poWJxXFI
YYfO+0kSg2+XSY82AZrMV3jWjHRunX+xPitES5KoGVjo3gNfE+JDPApLwMg7UbCdduZV0mvX/kBj
n+/VBhqCyJXj01eyTWdd+qKh1uDmUOXtZtUX8C4bs3nZIdV27KSV3MscUm7ewqT1m0N8MPGZJmSp
8Q01LjJzLrXY0ymfEn1pnsE+p9dfCWRA1UQaNvNrJ9FsWCU1e7Cl3qQjOlqZnr5jqSGrDeSgSesi
IaKH8CgbU+BlXbEQY8hY4JhcDjlfh6TrtRB4yUI2L9DglLx+K9YlWQBK61HZm8treATNkzbhMp6w
WpTlXyAd5AuVTfgb1aXQqdOR3uC1Kq2i43Nt8XNJTL/DrhmA3hDVWr3TjoiZktlGC8YKXzd5vtLw
NiZ92TL7XYCRJTJNi1S9Si7xk6i0BcW9gN2ZWcH4XvtxlurijdGoTtSolooUgZG4D/++9/YwnCCf
siyLkjaH2KXO+al25HVYIJu+nV8aogLFy0nW1q57Wt7KIN42Cp/come0v8xkhuxfCZ7iscNaOAyU
F23XyMmTxJayCIBm0whG/IRdIxOcFMqOhowvhiqe+Vznabonr5rkgygE5tAwlmctNkkR0uJNjqU6
kuTsYU3QY7jZs0v6nt0mC5mdcSFYX3Ke8XAsxe/cQLaVa1id0cmQ9CRQNS7U7Su8gfdrGodP/wt1
FPR5L+UPCGJlgTS3OBPA9KDIq4X2vqPbNMkZCqrILfWXIwJe4kQC5isbKSY3+liq/iMk1RVWBJ/a
UnttjjCwvOYkAOXcEn+7GQwwgRBb18o22gUfSBdgzimv2RiTXUKNNLSDB2fhMfHwWu/JCCnTPcyv
BnP2U5IoMZJRazWVxyq7DiBpvPuajLZlKuUoHSi3B5pmucJZe2z9+mPFXYYJtQAvYPYWkc9GBoQ2
+FXfn7WGRH1dlAdaX00lT8SkXgjkS4lBj9Rq+sCsUgiOy9zsIPdpXfGq/0yClVD2w1IogD4+4k4u
8ZaPMwUpVmaS+PFoTdVnOw935sxAxlQ01wx4Ynfq2LwcMxDiocYeYW2RT95g5k+/4eNKcdiXyKdM
w3stDyN2jf9ug1NrHxRy6tMywhre8ZiIt3DZ5ccxWDG83w0xesyG7asCRr+L49Xe82eJqdsmd/x9
SOJyQGO21nqlKIQ/fJcGj9EP8orQavDUsy/OJCAr19kWOrZr/13Wj5r/edFzXLP70rLPbUGs5eCi
BzmAkvJf7tZQEcrHQbyaUlDdjbwC9tL4wyxkcQZkUH9vtNT5rYwrN0EaDs1/OEbzaX6uCrMFquep
DAyEfa9zBzMnDt2+aJzl5KS/YRFNinuv4/zw1eqYhDilum6Vr/R3qSXEiM8UUgiupPUuZBlMYjkj
lQCwoYizhijZs2L/zXJ2NcFCeLPeqD2wf+IXpiD6q1qPn+FvRAxB9HRqsiiwRnRYObA3fEmyMoDb
aRjsRfgpLNdlARfjbTsUgB/h1+ADuC7F/RWuqq20LOU0PvidF4PWGG+GDLb7CS94I9dHQmgmYI01
UHFirVS/oLkXaC9mzzkTM/o7x+wk0J2Eed5x1Bwk0Rblw0rejVHidY3BFYI1bOtSEEmGCo7z//3b
A5VUBWTGyf13vb0hfg4KnVpNOxJBKTfQGMK+/lg2+SOi9CSIMoqaY5ems9Rd7Q3FhYThi77J5+nu
NAKj73ZJHQu8otGETCj1LTuSOZ4TKFeHzipvK87hAdbRU3NPvZuAC0ShJ8rKG9TNnllxsCgE1Ypc
CIaeg3R4zg/m22ALvQy1MClLAkFKokl6iAc4DXjWrtpbLdE7Ok1gcCHvrCpX4uF12ZbAqxBufGsb
Qgq3QJg7U8GGRaV0bgmftTxKODoZQNK49zRd+JPr49wVFjXuTMgWlXhrPyOEy6f0+ID3625PKDwL
nFngsSZH6e5vw02vN9y99sIW2d7bSYC9BuSVfBs38F5dT6grKaYxm52QqusHkvAZzfDq36CF8eC4
EiBscUk4UAbJYXColL4oE5+Et5r11qeF+k1EnbuuqT9YReBgMroRYiEfZs6wJ8dr8v5i567WnQKM
WkQvfHfDjh08jPXi2i3H+vx9XZ7bmUkjDY1u9YCaeYfKxNsOaHS7UfIaRmlp5J94z8ZY6Yrc3JLw
xMqhimqWBDIlaYVzF1NaOxndhBqcO+M72GYh5KKOnMi2Nh+qykdPKqZRCxr592QCDE1QVrFeXp3H
EmU0UFmiEzH3g1DA1gkIv/uzAG7/aJKnn0j2kR6as3Kjfjzt+46FZAy+xc8NMKlRvyMNklGzpX/r
Boe2vvhziufT4VOahOpiVEFpO+BVjPPNhfsQjpdyatcYDVJY111zNa1vggbCiwpNJPqOCgQbCizR
iRu3fbSAZSPYmV3hM8QXXsb6ZboEjpv0PyPTMDlBXFrJHiNwwY88/GTQMfXCVmOSoeBVFdb4fANm
KCr815Qmxcn7JmtSvBRCO45vcU7DtYpd/3KMGcvt2OC57N3XcSVEHQxckAvDf5lj+arC/7gIwwBc
53GEuog3jY6biq5KdjjGGcQpaRwvjSrnNkIYEHrgw2dqzt/uZjcsd9gDsX3tqfTO/mShJC4BEaLz
QBP+RQRL+AaX7OxnYB0ykt5QAMGp4+HNBtVRbrhPRwA08wFeGpK4Chpr3Y8n2MKlMFhfLfRbovDR
qNpZc/KtQvuKXUxDC2j+k/Qlu+eWBn6CUl27Q+jyyh/v/l2FGQDd80+8h8n40pxMvxM/VsvHR45U
JEs0s93pY9BHBGlmSc2Sk4aK/CmomgO3tE5ZnCqKNuPW5zyzttQtBWIPJ58PmLcqrmRLeEoBRlVE
/eW0dAmvKQlR3ucfl6GysAZAQN+kKV3C1zxEQGoS71v1wk8xzkSeVcJsokqrJcdabqgQXmlCU5U/
fpt+srhO4zfs4yyKXQ45C4kuHXabviotRQprqUpwWtwwc4f1H/MhVW79tScKGbNN32WzZiDTuBWN
uvlZlMF0D0hgPBk6+1na5VB7y6NC5hZyaGvT21EM0WErDSMPp0qAzryfT4Gp1vBvdc9mNRBWSTz8
85XJtmL+f8RHHcygaVahzrMTm7J0gwtn03ZtKs7jr/2ZbI6vq5dccYd24R+apSRJkmwypE6uubbi
0/TQpLKWa1Vn9cyi6AkwdQviZkAJ7RcVXnQLR2YC+67nFpSq8Y/eK3LBaR8q9aFjlgvrPrn/865D
E84Uyll7FtN8zaoHx0+YMNZCyPiVPRUwwxbGkxueLncauvljHD5XrxEPsI6UMpvmTgfKWUfGYHTZ
cPK3BC6wbKezfLDd5E65eYw4V4ol4+cRbg5+sDxLUJi3sB/F2u+VYLJZZA5EU/voT5Al42JUbU2z
5qiMAtANthXFuoGf6Y8E0uCMhwoDYfSWMQT+IYVn9ZOiOAlLoHHLBI1dVujVYAfkZFOG3ozCFoSG
Nt9Sji3mYViHdI95tX7pBV46R1bb9U/aOMbSCo92ACVV1NdPZYjKCItx2Gg4+KQLiA6omsa15CWY
1IVy4fcdlcsp4pusnSL0GiuvqFNavleRo3mQLnHcuoDC957PfHFzdBExwUcCgJJ3pVLIKebb/PV+
qAzcnrQ4cNK3SRjkWqzjSuB7o0/6Frkps4xra8k1fKGitySLDYRv3+bOf4KZXbC/vaeocYWgzgDm
ywFSuXDDxxmsH/pkZRYn7eYjB8z05mFX1j7KIed5c2RzCCDyFOaTNVFBLAGdAawelrY+ETa7N5O9
VGEZAM2zBAvLhybhRD2lVlIJjyMe88/TnWdCjvfb3FxKfPyY5TdPWNuEUujHIYsAisHDJgyKIIoy
ChcMn+9svNIiQHTf7HPKXKpns7CMZu+Ygfw/rhwdieE1fpfL0aTMHdrL1wVpv/G41LMKeG/5sL0X
d4PWAB+enwZ35i97MROb2xmLyMoeIn67xmEVcryktHJKsF/1wYbNZk8thwA2qsCC5gAbijnsMEGK
WLyS6pmTK/GnsvuP9D/CQl/v9lzLXOlh9f1uizRexyGsn9q2SS/sHaFh1evFkWYu5Cz+S7BJlQ0P
g1c3385fUl7Geh9SJ2CqUJegt88fYKsbNY/UuSBndycGBzTrYaLg5xEd/y2B6tio/TijPfmAkIwA
YHW62JLQEFp1VBZEYzO0NoogMgAa+kXwz1F6KljM5fVYZ7FcC8aHTv+mUqAmKe6FqDD89aTYoGy/
AzTPwfjS0YqME9V7AgS/pyTt3y6SR6eoeEOmGdqw1Q9fDrOfITtQjlbJGdxeugAL4YcAZNy0ZXv5
vptgU8aNdwuC5PCw3lqJs+nAaO3SxtuEwZ3D9kUPVU5oyu8gNlcbPXypMmFw87FUoZAThu1biC/0
EUZvbEDEUgJniGOp24riyR5DU5De94O1kf5eDP0F8rd6GD6oynULppSxdYc2DTytAY0+H2PnYtnz
vMy/QhX6msrw6jTeWYCdlkjkg1/YdYoCabPRYH0vtkZneKVDnbAz2op2p2iWg+ixTcaJo0VROcLt
4W5zHga6jpG7x2/L8DUoDeB/18pjCQgxb0oN2bl+X8j7imJnt7P8lcmPN9QCWlzWAVkMEk8dzTOK
BOxSJ2EuLDkCgtPSu8xl46+vjtpm7T7QxkOt3JJkAkvM605vB2OVeWetFsEW+E3dSJv2XSnJ4+SQ
sJskjOBcrV0Xny2eqQsst7M7v5ucusk6kRRGVUrt7XyhaaiV1rWxsLGmTjHxSZfYzUAlIitCA+FD
xUO4VO8/nCGZbSai/MjKniVLJpBxSPxFbvi/BOQKI3c79Jm7tWuAhqe0k93opBv2XHwV94VUc9pd
YHIOVNqzyFsYO2f8TzPq4o17YPUQ668JU+g1uCrqjx56GZkOYvjFGRaQZMPXR/xp1Knv/23pMEpJ
gIz9FqLZHJ1OD2fCMAO8+FseYyHOwGNU8n4CFrJMT3DDFBFRqo++v1qXee4Fe5TC80xNtAktrk+1
WK4hlGp7HusdIaNWZ5O3VthEZASqZ+yYV8hrD3+TA0lLOwDUpumvdtiH4sbyDBsZqkO8SQEbS7c8
gsqbU/ZSioDgS9b5oVDzr3+n4ZbXjLQAswVkmsXWeY8ExgWxnazEVSoaGt/94tHn1ixJgdcuHPd5
HnCMbqrBxBDTMLm+uskfzz2QL0ecn5dutkQYWmomPaTswaGct6oyz2wBiDGxq7+r8WFFvYhrVB5V
iWuALQLgYnbSsLrh0u+BzcoCVjf3U3wTXluSR2ufBOEIsD7UzGrX+d+TzjvanFPyarwLm1p567Qx
c2sCfrfRd8yfoH3AaV3uixJ94CEqReNqss8/DDvn4ysMxg3cFxvw7289RtnrYpwwEb4V7SPgdFUD
naUz61VKXThODs+gd5bkk0C9lR+xAL9nipWGEADmKZssmBiMcsDb98HEf+WF+MGRqByNU06EuaME
9RoCewtpAdKLF/bAy8YeF9siOALWrGeJdbuGBC8EgAbiL02yM3ivedihOqMgp1/ZlipG9MuoF3U8
7XSNa/Oo27kbE0yPT1d/aUFnXEuZRJl84fdkHILvPGdie/4aPHzHlHAEw6fbCAZKlWYQnjUgU5q8
B4ZLnlBbp1zLNIv5/aOHU4scxkDPmSPJaNEcyLZNUtrmkge0WHXOqhS6NsiUgDqZHU0pmF+gEyfu
GFPLLHZC2Kah8FPiPtvF8MXZA+o9InVfGkp5i5zz/ih81CzNk1zXhyZqs96M0woXzjiIbXOORhcr
xYIsVCATNJ4YgB5zfwZ5zWxLok4gExi+tRIjCnnmabkOmOfDlp6sdfk7AHcyR7txEugsstFb2X2k
PRcwG/EC/qi1YtOT11CtQsBgd31C5XBVk+mM8Ro2ruixesPQ283qzO3DX6tfZeL3LGPQxXQuMK21
dz+cKnBMmLvo+Nb1HtTct39n0E6qPUUy7y/+nM4uuZlVAC/cng/1IXWokrl4plHjA0qL0W4VY3bD
VMDdEFBcClOBE/c3zV9REyY2xeVjG5VU0pdjUg1rjTxGvoYngsSY3JFdLNENVAQ+FrVpA4dP2m5T
I802KaJ5ds/uSS6PMlt3v12J5TMzM+WL/LxtDpLNJfSsM+ocjCJRPc4IkkcI7XHYFCYibNKRZB1d
LMrR8Gt5/0mvjFwMXyYDf9tGl5uZlP6YnGMq+8dFS6zuO57q8TkoFVkVKCGMnPbBItI0C2TkXalP
sKShSk7Yr3+zETF4dC7wA1c5P+MSHZiMbO9LIzXtx2avxpEth79vUWEiv8ugxUa8yXQ752SPPCtZ
7RoeSMlNV9tjdt+I1v1KqzsDaZvVJ6ZdFUelBwFHHCaGthV/fD4qHZPBPbgpEbezmPqEp3Fp8QkL
4zuTqLl/0gXRqnJJ/pt39dwC7zKbMEzS3jFNwYSTUpJhEK/SrOeMZd218EvbTa5V+b1u9K2DddXr
1L6aSH0LBbADeUyzASEXJBG7SmFjqgXsJzWnMCMZF53A5RfM/FhytjlCsrSCCw16Z3ZKMOsEnfeR
FLd8fTWTztl6NvHsgh/fFykD+66E1EmToqXP3QovFPo5GOy5uI8kPCeahnL/szLsDM83o4/K0F70
gHyuBifaPjgNa06cgepYLFr56d7qsT77ndNbKUdOEE1f6dXwfnWJm8TAC+90X3PJCuZuXxnQeR3H
Ui3VYtN490eQP9wxde4RVsmZcnmWLFd5eDSrtgRaSpDuouU9ZvG5Tbnri0LVxP9Km+AgiRcwLhdc
uwOsv5msnMI355eXZQL98oVZ+LRrHTcLQuKII6Z6wG/DgWlFsZVyKQzBGPomdI2RVBjS+JW2Dl+I
oCxv8dUZM4+S/y1xgPbgjoJQmlMET4t3NjD0L3GLPecpyPFPfRuQtJgRiXUYe9BgP/kidlhQu8e7
cg30e3l1Xq8lU/UPFtImyCkHj3a2eATg9ylgtHpAhQhZtsCM/evR/GEECaAHoWO7siXl+4+dQY0H
WfFrrqlJNL4nFolwJXzvCuMgTHMZuLNJfz17c2p1siTcf0/T7shDTO43nWAwerRMkjZ/mkEEvtRB
QmuZx9syf6E7r6TDjSaEV6R/E36twIkAigH/3scFRlLJ0g+A3dHyoEyvph84WPxszmtVjIDyhu+J
Obzoq+mV29Lt8/dpguAaua5ZI+nV8Mt4uCfQUnhdVfq0hNbInXQ1tsKaANH8jxKzbXGlroh2Lv4w
XAQVGZ7GeQcEWmW9uzZbeDccYnqGf+TYsjgwvV2K+3I1i0M7dsqSpbNC1WjSYK8BT9215eBPavqv
Thx+bKgNWT916Oz7o0soSgY74/uLWPc8Ix6sJdljP02JSQd+r5plrjJHn7MCGw4uKC9NJBkBYrZG
1HIdLxk0Dim6IMgFRUAFKGRXvfDCfzTtjtSMm94hjPci91Ms/ig/qttMKF1NU6fj1AmlqyXKr8GF
PFzNkBGNImTqE7RpOzNhcrOao16G+V38K7gepiAYOtBeMl1/ivkP1aNU4fUzToQcenT8ygdixRTA
JS1WfhjTdJZXpYmvaUcEzY8B6GLvmBgvrmPObROuiaqJkKK1UDj4gvEF1cwWiCfp/wpsjUodXZPl
Elt481R2P/rR0aoza4qIdzovR6ijNRmh436Etikdbe5LHI/QbV1ywJ/rer0gcfz+0qQiwgXT67lq
FxCzcohcHensQeKlaYB5jdw3ZfTKL4LBhJrZXQomN9fjxGSH+uTcGJpmAkGnSRbbAUPi1LPaMG9N
WceCa3dFqTV9YwPIeHxOdhdBisnXPrUrACkan20vzMOGUdMw9YbhiXHOTVQcPJrV7I2c7iwFWp7T
suWhC8zPiysAjIIQrkzTLoahWdDBSG61UHVxmycBQ4eBKsfjhsy5D+OJLSXlwxqgsWRfMFvGOp7p
keoDope5cDv6nHsMiKpVDTkFLveQrA5NtxNzOoX+Q1dHmswJPKZ18RWjM0GgdKjcvCSd/W0KoPDY
fEz65dmMwBEJfVhfSAY3FrAnc4HBcp2Ilgf9hoI2A9Kdnc9SMMDHWl3Do2dw2GjaUkIcSC8DDw5+
dumCM6IBsDLxUStmJty8aU3LMYYoREQuXNYGZj64UPlsilcZtPSrKBxxn7PrAgq1aWR1vZrGpk/i
Tl79sHJ2gbE0sz0WoUs/EPMSmvw3H0Q6wDJNdekk3kVM4TsbaBxGVbaUfRBQDO8hstEsdTEaUWVl
xoBPMwkDVED5bT3+D2QX08Z26SvKx6cQlhlK83ZWob0dIzTEBf88/OHbH5gw3eEO9y5G5D0gI/Dm
4DGRdfRTOAAwmDvoobzQkQQQdF7d4aIz3WR3l9K/7e7CC2g/dDqSfAkJPWfQbQvsAdWTNvs3LoD6
4i3YzXAuixORpoFZxWwcEzILI65OQBMCDnlpcH5uokWpkCkcLCnWg1DP/Z88cPYmmK7EKUMFGGLg
AUa6MPMRgq88b+kfsjnQQK8lFNIU/PnzzSMaQc5jAlVJAC9OVm00a1ubNj1DFzssEkugcoQA0NL/
T4t5eUMxdvPRdF4I1XeAa/hGjuYFObq6I8L5K8WwvGhJQENZE7K2LwF53RTJH1SOZQBWOg5Qk+Lq
nxWiDdd8JBBH1YbT+LTZwmFIza56lJn1rxY8k22Nt2ttJC0a1ABudHA1LYzlAAIIokjLa3672CNa
9dIGSD+2qCdeYrdY2XA5GqqY2iq5tPD4iaEiU04i5COYirGPJWVUDSI3NWANYDvM8bi8vfvSp+hC
ZoKEkeHEdWzO8JQRcVkLecaAe3WMATQxwn3Dwy7qRqnoYu44FWUA6MeUxB4fSvh5hFLzvD5vNtLu
cl9k+IIf+/xRlWCbrV17wkzM6Y06DMKvuj64x6khZWf0AeZ71LQPuuljPXBosX46S8s//hP/49bJ
3Zii2HKKBjDd4eud0bjh6x/HyohmHtuplJoXYFOol+WqeaT8AJbk0MfXbw904cNajNCoTvsiUrGi
3hOD+svdt94fSTjXUqxot1PdqiE8IJNAYeANOjlTiyCy8T4oE6YXqegWwNXsH/AC7CIFfrPk4YSe
XOKc8oxYkrzhQmR0fzfC3rqTLfwQRL8f29xb2z33MM3e5KJAVScKnx/tk1Yv8wbHCup/tkSHuIJ9
PrpTmoqP28FlUbbWnP+2yw8thd9j53MA5dEmD/nymuo9e0zZDUm0pFpt4N85HErEGXQ649gOqkKv
nCiUfFe/gPFwezdtFWptxM7DZbor4xjPqaxciapg64yYV1hE9KrPYq63M2i1FEvnWC2Nc+MYH24N
obf64s3ugWoMxHUXtI7v4fCVM6T0FPdiElCRHuVoECOeBHERb6Cy42qaR+vetpfEq1zFE5QZ8nxD
+ZwW9mLxkRlfns7ge/JoR76lazl7NJCvUFhTD0mNTcsaw7kZqnDv41xPt3NYxK0sEsaBi7170+1F
JiF0z++OZ77t3sbDxDUh0ZmGfpakx8EkDYBcadu6y5uICz9qtfEARxwiFb9aSjVUF6f+o2tVE8Ag
8SjAJMY5v2Mxx3kqBN+ayezmSNEVywgTQIw0XVgOOoXTXPUvi1r6rMVvCCKRaa9+cSeqcp79Qqcx
PmsyclmpF8sl0e5fkBvX3jw2YhBfXPG3OMPlT97RPyDig3ryv7zE0Ih0+INAGmZHvvArfgsugpvS
BuL3Poc2PD9CaDVk64cX7BY+0lVZeTrel9lqfH87ceFmuvQXNKJCctvbmmgSMCNVrfnwEdimycD+
pfgB+U2ZvBBC46VBY/LsNkIbIhnzY3FxTw/VML2gVMWpgS80PGak+/+8QqwjMrsgW1tBrE4vkDdw
9dQGrBtOrFKPcEtLXiWmP3ZQfQNsSIQCFYPqspOLVYIZPI/LM6tKOoGij4r/AxWHa31KoLPFa7f+
Sm5xEg5pD/AuUr5++hGt6AOI306h+0DC7oNLLOcZcjBGelQWhlvcv91pOFWZOPg/7D8yXGob8aB1
muh+jwIEJkzOqg4L5eSjd3tQdb58m1+y+/q/ygnIqyWzCbqpMzGWSAOVYL1Oy71xfWBCfF2AbBqe
KnGEu3BJm4gX0XFjQXmy8JkDgLFio+8wjcy0RD5vVGEADPBeTTxZGRzRLSWQL9Q0z0J6iWZ0WyeS
/9LjKcJ4EWYWUxlY+xrFrAbsT41QA6ew8Fjrra07S2Hq46GXCBUeshi+Lcdyr3DAZ9l1xwUkmrSK
AUhUN8jvTGzs/uiHNx7KMytDBxSsMqNDGb1942ih68kAzQimvqwyafk45tSmP06zweugC4joDlnb
A7WaXNgmZN3tKRg5wut6/5NYxpFIJuMfhulcjEwGVuK57MAzBDF2wRheHycFRVu3NXAsR3D8xB7B
RGUewdmcmMfiftsSA1x4EjO/7iUv76NzDKD6+qGBhjwFbSxHJ1NDG8MLL5wcpWunwXzA0a1G1gJV
U/KKtvB6zeTCtfvSh3JQreeFY6pX6euzHnMX9p8kwEyEsCBvyfgdmiAuUV12/hundPR06++hwz/g
FhAHxAU1clTHIKmJ5z4ZMCCYZdJEjKn7ElfkRI5kv1v5m0TRFcjbo5Ut2dW95hd9XpswodVlH+zc
5JrS4xmeRKD1NAbQz6BC78ZKtaTdMS9ih9/sBdRgC6AeBNfC51R4ta4yiv1iaYoWy64eHv2HP6tE
HgDv58+LekUj5UP2vf94quqg57et/qW1vFKgHi/qeN2r5hXMOfWPcHxFtcM4GHM97TZuy2lKaKbN
MnNvqEF90iECMNvLr4KSp8Lv24xd0UWl9FJHiq6zvyMo4YubeeuO6j1iJxddLffSq+2M1o5ChHng
imfLhS9xrddi26IAt8H3EU9wmfFA1Q6jxyDYmvwmKSyHeKXq6Q/cHRruATWLZdC3CEDRKOjlfZk8
vU5ZVNhBma8bmntLicSWGlg6FVVW40PltYWKPyDboXQVGXQuMGeUoUCMWbpnHS8UpSbHIxA7YaSn
0vvvE30i3mkSvdX8w/OFPUVc4V79iydaiFIcKYaLTCKBZ0Zo8EDeNyhJ8RWGgXf0Ii+aJiruQrKZ
7LtjYIPISxtJeImelOY7szPFiAN+sYWGcF3fteOT/OOBEtf4qHBCE1l9izslCLmLYNOqNbsc7WAU
Bpr62eiQEQDLpX4KKtQZENxEhA8Zhjcr0Dr/bmm7GvDWf6YYIt4EEmqa7jpqIRmf2LAJhB9IgWuM
dMOQ4W133lmALO2dXg4h26+c5wIIJhiX7TwQDFevpB7SdIS7QUK11meamdFhnc54jCW6SbYoATy1
frph+LfdmY8ACvuejAoius9Ez/5S85ilI4tpfPs4hPJLe6KggkYiyI+lbnGsJP78Lap7qlYvXefv
pe2+TiY670rIiYmBG4senPmZcPfj7tIJY1zcyWGoB+7hdjkcTdtT9St6R4e83mLTVGMagzr8JjZh
ojx29tjMzDy6PrnMeIbSk/FHLYtCg+NQaptelGRyWSO5x/ssG0GvmwuRcxJ43BjG7bdiuZcFFcMz
w0Re2oA/I1Hw03QcKcPgAJb23s6POkQ8Nj0rxQwoVlCi+TvP12wv3D00b3avOMdYfwb9n2Dplw69
2cNCPFyS5THk1mHmsdPMCCM5ABCzZIjcW+PreVGBvrNDwnHJIUcGeLUZxTj3PWOjQjUs4Q9Cpkis
vcRGhPrWs3H2tguZMHV9CXyoQ5ESTEtPd+A94fbzDZEFrCMhgSwLe396afzO1P8ephsGcSctqxwj
kaZlIL76Euo83kdAqGWDuYAe2yGCdT5q8egtOOl2OfE0K9EBhKNx2Sv146YRqgdYNxZVHVjDCD8G
NP0+1XcPnwHk3MKjLyVPx5BjvpHjAcAZ442QK8pAqhu9hAFmGgoFNcdMoJIrBUMY5RG8SUB6i+RQ
gRMPNPXvB05OzIMoSnWFDesKKXYuWvl59VFfOrW2d58kNYUYXCh61ZXc6vd8Bk6mFLKd010wxKRz
oomsKzfKBe+ZmIQzfFP+CYkl6DO9RvEgjFVKsEdEkWIMg08nXVeadN8U7I5QW4dwewmoQlKxhYMP
OUwxR3/wKx5LkIN5iwnimKttoO5t2geMiQLeu1q8UhFB7uEAm+Fh2PD7cbD0x7GPFF2q8ZtKz+Ir
TUXZIth53rEis0uH8oHxzMeOjQP64tG8wkPl6ARxae4I68TnZdkH3LgDNSQRr47q4TThUZG8fLu4
zrEZlAu83VwQDloUIjUy4IZXr8f+cGkXRhlatsrRh/uYZ6zuIGy0dBUis+welpjnWwhNLs4k2BPd
eksgHwL2LLpTi864z0RRy9kDqnE8aE3vFrMws/ymp0dHzMqBBTJuLFCBzZqDCTEQxe+Aiha+cNKH
LEdQ3IjxKzI/xH/gqso56slMmiojSJycd5axOx6zKGRxZJfLnNC46fHXk2Qft3lYFtPvRf2ttUrN
4APb4oveiCE2jmmZ7GMf+S2KhYcIYXNWH8yRWv2F5+CnGbhHgrBG8LO1W7feXIbFuRQ5m/3f6myT
2WaP+4leNtssCW2JUm7INbk+CEg54XOO4tJESswH4JkVvt+v1GdIg9Lve4cbRcr4+RMYveXBY3UR
qTphPNC16o4YE8BRpa7jqZ6dtoJtmtRNEMHNih/V+EEqWuQsbOUovtAMQJensk7RsUG9G5315qe7
H7dl3Vc3rrHikzfLt6oE/uOx/M38iVtgA84ryaXNcnZ+U8eG7JxkYUrtmvrCS+sfzs7bSG/sLS3F
s1T4KYUe4f6isPoIJLGvnfgCKnLAXgXWKzveRHMTh4yeCQqqPrwJiptqazAHoAFtrr6CzNJxLD6f
bncTHO0BkI3MKHqY371DVIsVoblnUhlNnSAcFef88IP2NFnyfVLslbLTDxiDKl0YxKrIyOeSdYfi
KASyskkUor+QvshnIR7UfbPGQLDcpiB5C0Ez1paoJVWSFacJlN7ueISY1VwXr7TevwhPYiVopEda
ZuFrFNeogYhxBR8GWdK/CVvgNaYjDQVOtlwqdRuJThMHbN1qPzPnmba0TLNn3NcDUZ8CZA8PEPTT
LVbjg4LFo+iBEI2/un0T1cT6YmfKXnxT/G5n/tZ5SiNIfV7Iz1Q8GBqTWo3CmdhKt+KDfYb1ceu5
lArWhimrXAhERydSfc5cz8HjfTef/XPUVHOyBr+9714VBeKfXjbndMb0cBoOHhrrvY7DctkE2Exq
jv+MirsFLoGeF5vn2Au1oPnc5YoQ1EyG8pHIRDtmZ4n8KygpNAb5hAdgKun9zo4mT+RsKo59bQqL
Y/5hPAoCnytnl71/AADr5UAQE8TXa/sx/fsI6gGcPW6PmOfK5T7gBmoLx9M2CnjtDP2XaZmiwF1V
nf2wJBYNF69kIhQACKu8xTTfM9tFLS/vjgI0/N70J/VLBiKILYVzqgnsyJmX1daiE9JagnTZlnjY
odFxTHdChVCqj+C/tY5Gmbkp9YfL6Obu9VnACJBbEa27NB+sRPde1tuDy/3n6X0yt3pS/UvkE+7Q
rr4HD0Oa4j+wJuuhr5I9H8yGgFMUY2sh7ShAh3AJCLRIXYitrZn1OPBNw1ndG0Iht0CpAqx3xca6
LnmORZA5rLK3ytck+A2nZO3j0RjpYs4QzoiMO6lQlDxFHxZHf4X3P7Kjrb0JMCdwBZrLIW66fzWt
eor4Srb9boAjaiZLJWNBzXJhVQL6dRsq+FpUnHs1vr3FcJ7sB3/sx8si1iTKyNJ1GVPjiskhTqsq
Cvx0db7+tMqIfbAsVZkz/qJ15a9P6Fll7525OczyBgoURfGREG5f/0SwAhidooqAhFKGTFTG7mRw
GZ0S01mqAipWAxRGvH1hXTYyWGVh9JdgkoKHMfVn1SolkGxARuL5GzjNFLqa1GHPDgHvkv1Vs6PO
dRywuuE4+cMnzLIY3QOizmEhoGdSE000jEu4xB24xlot8ZU82wYfBMASJUXX+hh3ATkEzObu4J1X
el9i+fvSD2YQ0KiK+JT/NJk9g3UU84NqFmBkMKjfhFtA/g//mFMDq012eDL9OtdaYywGU+gh5h0p
gNRzj1jL0clsO9Of2iCVM6Kh5ntqkm2IaCNlgrOhGT49aFGukl664pHxzxyTNaGCSb1Y0mHazVkY
j/hBln4KPZS7kJHpZTxJdT2/9N2nA98OosQ2M7ALzzWlC5RmzPCxLXuZrmrf+2ogVNdMmxQ9aTk4
os8LBU90BvaYGlTzIP/jJAENJkUNzqD5O/zagi9mx8qbxMaT69DAYDnQOSKjmTJVfGfYGEK/FZah
a2CS8GsymY6NSK4BwtDaHGX5kmvnox4X7mBnQeKE2oZu+0Ez1dw8PW55hIagZDsDSUETikvvFMnq
lEtdXgth6oryRADB/VwMTO968dcQ53iQu0Xeu0sXvodP/eq8U+4AgJ6TcQlqfeCNv/3QEkdB00xQ
mCIMsaMxJtPFCcz7+2JNR4Ztt06GxQO7kGLSY8R+33nk0GyphprXHljrr37Lze26vcbmZd2/Kr0J
sMsBW5aVdJc0BX+Owoar8QX38WJPowyDE6U/vkXbzP5Jj1bKo1mTcVhTp0LrEwT8rzPg+Cs49VRi
GuVP8UsDaAQRVanlSEdbqkpwKhJgUpM6+0skmz8uR+K900l8/GvfaKKmxNVXfbqdYkzUwNP3a1lr
IF35RdW5Ni3KqBYzaabLae2FX6GyIVv30CQinOXRuwJetx72f20wczRQ0xwj5l/eKdvl7H/kWU8p
l/02caxKx+NdqrO3lF8kSxZ5qQjKYxZOw1D9aFgYoGl0yePlxHD0lTUN7VXFeZJNik91KjTrJqtv
oBq+nZQbzBK/f4lZgbTaQuNyB5Jz0yngEMTe4ObYaubefRkXQO1tbUwatnRKs+FpXnlVs21oHpdO
TXX+llyigyjU6IOXM0R7WSMa22zxx/XHSFrUckNrarrSPEadZWJDw2NB+WtuIySWfcNkyXJ7TAYC
0eYGb0UU73Zu6yjQwscaVr++Mvh9kFHSuIsOUzaDiTxWooLfn6Jhz8g+M66YuuoPYErRSdbE5Ljn
KGNCbjdpkkhyWgNCsg5reZrWFjZ2lKUz2fyoYLvpOiacqda14v2juJ07rMIU6DNmqJhAS3RIG4f6
tGAdrkAIjESzOL9mukDO/bbTDkgY1dhR2EFIQiGXokxdFaXdhBcZWbpSL33KKPmWW/868ORUFsFy
0lJEN2yLMBfDlGyxwJTkpB4DKeI6D64WzGW7WnAsd5dNhpkVE1dl06dYTYXhPOdhjFNPKKvM6H2A
+ENdWwgCBDN/9WXg6u4cce5Z6qTy97Eb8TusYdyc5nBrnDOHZ47qRdZ33lXhHjxjRxYHEsVM02uP
2FrWB3MYEeGBMCzODfnkqkzgfar+6+GOgl7iMpK45helwicnCeZVB0ed8uyQP/I9IsTfopDy3kzQ
gNW1gB31BddkdBXkgtGyKTGcKWKuYJJ6pQexENr0y9tMEKpErfW1snZYIPvYuiLv0vg3NNlHT3mq
VpD6usiWzeLTmKOOf5t9Yq8QOzyqUpAnl1GZh63NlUB9BSqhRYju7UNPeW5FNtJ3n1gy47qBBVF+
NPl7vvRx3bHgGiHsz9Vomgszg5CPixU9Lti9Z70OVaTuwDlC5DJLPtmdbfs6ldAOUkDGhxnjTQhT
dOvAjy8I4egOwGspCM9OgVQaKAsP21ze0jTjaeE5S6Y0SIbJeqljziDwFEr+EroSKR/zH/L2tOUK
Jvo7YJDxlV2wTzSzhrY9yyyG4e11vNzXdzDmo4MDgJTsiCTBRimMs22jEt2fHZiyptDoJghNaayQ
g0QmPl8cNskJcFd0E/gdJ/ryRZCfSa1PItSIDEd9gwBYARyaLsrvI+gRPMVm2oe2wYn9+qk9Y8m2
4YXK4pW56HK0hm+EXVmZyoHy5pb7WfGDrsOqkHc2/zrj99ppWJ8KODI3DqkTB3RWrXK+7bpQSnXm
VqzRUiXmmlIL8eAkvG4WkuGMGbYOtROKj2t914znYAcZH/kH844GOLo4KPTF9Wc+xjnA+n4ZtXLJ
imXn70yo4P1BsiMC2hQZhXj4g7QvQQNjyhMddMbHIGGHkO5qfybEXdtlI7D5VSSeq50jh6DNXahD
z/irzUsUAuaTSXOILc38imidTcapsNVZ3Ws4zgh7Ge1PjWNIsZsHsOrgVaOlfcRCjUh05fZGfybN
QpwB/ShacCPMxFyed2AUrxT56ai7pVRBIoM8yXaJOULS9gM+Keary1VVYgVfSytPmyRVxHfwSY6P
VzLecU3B9LlhGUAHfrK5/lctw9ce5ApjoWfCS1i9X+LuU1OxL1ufDwG9Qu+A/zJ3x3k7VvkJh1Hv
Q8I8UqbL1PQu0qjKOKzAt/3Oex1UwxXU1+mQ+jvqmgMaSEQBxnzLd9khnv0v8QQyKvvygawgiLIo
ZPYuDh1G3tt/QUFtR1BCmq5pSqWg2zMrqBUS0q9HReV2BfTihPi1Q4ciRS1joXYPXlwDnF1391Yx
3GHHzNlAj52ZNux958gsN9wdnEc8koPajzpEq+T+fPCqlvYDE9x+PMtyxksgM3M4L4QUU54qNkU1
yluniuoC/LILPV5VHpY+haDlZv5S9xxO+6eZzt2KglpEb5S4n4Ysl7NMyq89h4cd10bwqqMfkY4k
Y6Lcj8jUncwOmjVpmHqYCU9qOeX362d5GeOBnFNDli3cKT5cuUUQRxIIScNnZYcPW3bomb1XAoQp
kpM6OYUnVFcLK7jGuelWLjESMiJ9JwD/pGNdi9y0vx9qDX69r29K+rOFrCCIRFGI/q0BmqMd1Ykw
470hiTUYajam+soSJwkia3AOEv4dhRIfjgS9CCe85HRspkv9XojVVSS32ZQWzFm4J1pvmH9auu7P
hjN8Bd8A5xL5uVJTLyFJOekxkn6u3W2W6BAZnY1pORryHHwyE1Z5SfybIa943MtQowlU8Q1auwLM
1LB55SpcSfgMOKei8BRpbfgsVZSt5X4DCRp+6rIzI4MgCdoNXzHyaDRqI86FCb2iH1KvUFxmA7As
ubWZlQT0bHf9ocshA/iSjw2ZS1QWIEnWCzlWaNbseDLIwzNHvuCFnh7CUFvxt2sfRjBEWvRQEfhM
+6gm5xUQwQEF8nqmqBkFuaL5yEDaDFH7MGT0GZb+Hov4DBu6f3nz/bd8NrGTt7pvpJ4UVKWhvQA+
RavPd5g8rkl3xYADl8AOSAcEpH/9L9LUs2kJo10I1/VccLqDeG9IgulDqsdMy/OrN/x5+U+hRgJw
dYMROfQnE8LyLE6lbWMRLJCuC//Xf8lc4raEq+kSEObj0VdBZi2Vokq0HJqRhetqoYpUVoTi9huA
HXpq6/lX+aRzIFfdGsE8s/flRrwXrDJBEpthx8Fq/WVw/JLPvIizO7Pa0RHkscirwJdgsDyZ04en
PjptUhffHG8MGTGeqGdosPNZJRToyZb5Yo1/0cWRp2p3AgnSHZa+coujnP63ltYmx4mKal2mWOb2
l9a/bYKsmWFhL1m0BqLJWDveXwIlommLDqZbhHtlAiDdLGrrtYdDa2jJPOav39zgnGRAHAAU6CuZ
ELM0hQxNO0iIuHVQ0PHZQNvAZekyqVtBXe0fDURRJAfj6Kv7Mpgd1srmKCdsTo1rhRycrP9gZwdf
/9s6SYfxa3z+cATFJ0Roa61a5AfjD5rLPS+YrDIo4Glu9gpcjTPkovEcX5d3KzTKZE/TRPBW0fUu
NosRO8O9GV3YG1FwxJ+8auCf8IKMAqot4wMlMAMAq1CnnWcOo7dx013dldLCXxA7J9/vhIqlMvdJ
/V54EDv14ERdI8hfopuBJMDGPhy7ObU9KDwQVBiY5Dcx6OvnR4gXS8pzh4NXYxx66gFaxGSNkpyD
qyQ5H4+G+VbGmLGUio7/GF+CtZjwsoblkd1AhSO/6s5GtwP1ZkHOJKq8hL34YDaenFi54MBsVVvi
ZK5CYwSXE+7bFPxgtJ4uccYqdf5wjhjXiGVgeUFT3ukn6QhelNSa/I9vOG4EC67ArS3ODyUDEPwM
tt4xU++rz57pPT+opXoNGza4n7j0IKkGBybBFL0rYYNyiM2ZsutJ6S+1soZ2c67/lbSwdm2GWzPW
fqZrd18Kp1PEuMm21s+IKJSipe4w9yCbay1zjQCM9EjLcVRJGJB3ubBH5yp0vzm2RKdJc27Iaa6n
kRIwD6s0+g2JAZYnuC5mVd8ayqWuYiScK1+kECIAZdbRoBVr8fncQT8IScGoJPNzhLHS1LhF4rV/
6wpayxm8UOQtReyJfqzrE5p7bVR30lZUKOPSCphdlrYmmar0LmLdXvJAOxltnhDn2N/F2EUXe8EJ
3bYqPWYyGdH5A7pVkkGN7K6qVTl1D/QYBmCQUQKJVMwrKB2aCkbd2yWqiZzxJMPEbENQHv9aXEMP
QthQW/QsUYZOItZakryClTlDqu6CzpGzK5NWQb3DipDn6HnNmICQZfhm10lAhbUHSEnC5KIpFdT9
2IsotKuDSxwEya0o8IsYV4gVs5QxWSDwqxZUN2k7nrFSyWXu44zMDlC056jt4WxrhjtpWS7wbkDG
rHC2Wsf3i4dbMabeXRopZOjBheqF9afbuf4AOO153Jm2m9faFxhgbU3KV2YOP1+MPFWAi64NZXGT
m10slEqjCFZ+RdU3ABtCvahX3ZD+/6JWbt08WpJOAzw2KNDn/uY+EUDEkwitWuTJaev6cIkQ5MBT
zE6VLOUUijEALz8OPArmyFjU+iifDTesCY5y+6jQ/oCFQPRdmJ3pLkDzcWiP9znzjWI5mf13mOpc
Hif1CJGoCec285EzA8hmwkPu5O5tLgfkjr/hUhCELgunW/KSmBfGogI/jGAhgfD6Vkx7mLVMFc4u
XfwzF9wUdTv1yRqMreKIjc4uoQxr1k+w9SF24BgdOnaewlaStlkWTxyFBdvObD3gy/Q414vVvcZR
HQmTSnAmfuXvBBRC+y9yyXfssTbNbY0vFq4aN3rkSXB9AuCxY8LfFWyOtAHxoES23fx5Lk+NY5RK
/o8uUpUKaFhQrK/gtd0SSLvjRe0uoEIDqB9fkcjwSIaU/3KPxLoz++mAwEdByWSRQC6xDWkI9wH8
3UheR/KIgubmV5YRvWgShApUBYiEFdH0c2QoZPtySux/aaQD83MRwWVmJk4o64udYym9NvxYeWfD
p9pVRnW2SKb7VNXDZvRW/LGFfYuOvCiuzY9md/sX6Vo3jkMh1tdVu85maLRQ/AQrb3GgFYHWfgjv
onj318jHa5HeVs4Ug6hkOCg3LMA/zqNWVi9vMw8BWHRNJqDaEr7DQx/yKcCx6ZKtV0tOS6+qGZO2
mmxSOlFg5iEbx1tWOZIWzGFAPlyJmL3lZwBZn5PWfiex4YS9KRBNMSrWPZJwYQoTfd9S1mCxjeQp
TwWODM58Ux5GcVjLrx/6CY5rv8Ww11ETNeSpUL7eTJ2jWYamR7crs3xyUBtvoLhVejsrYD2wN8Gx
eWUA4DFzP0pMtZPAi6SaSD6kDRF+eJ2xAi6WwxWO3JU3O0Hh+gpiGjojkKZC1VkQ46PHiJOSHRbR
mlQ1MzAHknX99eq/9SLCPpld5mbWo5G1tJs65z7pIh74CXG7V7IwMiR8mPcUZTzWqRCM305YupUS
KZKZ7dX3+KKpMCuCXharr8skNd1pMSUQyp72QE20eFrgbtlOcSisrk5u761wMK+4kK8+irAKLGMc
Fd+UyDO9oTFE9wnmsVB3uSwoXyqIK3GatHaEk8yffKD+GIifckXARSzl9oIGEYQS5rcRnEKJTu5E
AQCRV+/hYDh7C+yj8PpHBLTa5iIjJUzX9+8geAmci7SPweMzYO2UYMQfCZbFmUwoHPbrOkZ0fQZi
cERK8Fgpvd0/4QBMEiMBI8A4DLPHQMO0i4n9XdkFsb7wlDsoCrN5+fKfU9HEsz0DqADOpFZLchdL
tGHELRIhop5QlSfl/oeLBr8E6qLOnmLRZLse2wFRZ1pclUT+P956+9dtnorTRmMPDwSfBCohNxHu
Be/eaZkYhY1X5JMXG9igBOObIEH8mgGWIoJDkvx5r5XQzoUnMRm2wAeIHIi7BwWq5zGfBuQbZDuQ
nDu+fAsh2TKUKP+Zl/1M6IiEPsjD1RV1rKN6YDFtz8kANoA2RVyp2EGqzkvTW0DqEnlzi5xZDH0g
jqDVb5kXZZB8ZT/e/zMe/NSfyDd5HE1arGdkb6mwAjnatRMijLk1U3cAvmVC4xefbr+UBN5ukNmP
I0MSPsoefAoC/NbT2vu9h1ITdf0LDl/WhyUixoYhas+Bb+SupiKDlwxdKjbsax3epXGSPU0qMu8z
KHGNRzWlORlKIwEjRL0JTdVobTOg9WSqDGjerg1AbUiip1gVjq5+vlSxiegMNvy8Fry+FQU9qgAl
DQoh8U3WcgFQ7aIJEYQcZaHLFkPfX3FbXyQy9kjq1SlVIn+4D+/MrFK8neeFLwDDImrm0zi/SNZz
yYZaY+iPdIkjxGIDsPflXOUNUyYmlZI54PT523TPaRVyT/QAt0oSNM05sHgx9uh1+AfuSfskl04f
3aQXwy48SAn2FQgFiardPwR0i7V7nXF9/7sWwBnIiXUik6D3ecqa7+rOOLRRyGzLnYdt91hsM3Iu
9fnYc2I1ZvE16y6/nMavg28EOdo9IAhoWKAnm9VCEoJt2GUp2jYD5MyyJDPfzVcSYJltOHV0JNhf
o+Ys22UJzNnQu0Rhoc3/EvhXlHe53GTz/QWFPrePHc4b9FCw1QmCNgPFZE3i9tHjR+PXgrbcEhT9
zQl3kSVhG17Noc+Uf2B4/en/N6H0geIqzU7FeQDuAaFJmEPjIH8LSGH1G5g+yFS7vS9/Sb6KMUU8
/AXu+uOB9AKLWixNtXagqa5jBjcpmVXYsGmWwgkx4hD3D/586QMnwI9b3Cj7otqZ42EtvyZhObcJ
GOHCjpFXsiI7hnXrx9PS5vYlExpNspNiQH/RtPtjiKST+blcVjOBys2CNmcLOq7HuvMluU9eg5IE
tnfcXZLtlsk5HSHhBBbfM7vC/cVpubgLOmvCQNEXCYQbQPR9B/M6+vGqf62uTTknYhEsrESrOZXn
nbt0MY971sn0af4Q1Pgg/qDWiDfOuPO/kphZlWwCGTVZ0/aMYw2ZV17QKcfxCWhefAugdLQg2mTR
FpET+UJ3KcaL/2sG09gBxp20jGq9ky2Q9eUs74pKjF0yqpuy4XLUgJdioY7EpN1tbTDnt7idJOrq
6xbfWEiYxyyPD6H+ZZbc/+QY2WpSacxvRXSGNuFITlAHIGqPoTRdDrVYZygVH6X2yq3Bx9mnu6rJ
F5AaNwRWzNnGr+/JQKAGLa3AN8V3KunxT0V05dW2lpgdSly1/NXz+rw2TDoTLuAkqjW1nNqVZpGM
2Eb6hCYmLEN9plhzajS6izDgl28TIP85d5COU+jdpcGa7Q/J14toXuPP22Hwb+zebUSuDJj583M5
FUOXkXnnQ8qYvTRdE564goi2paLHvee1X8FNl+rtTnhS02ki5RM6rwQcnxDXPQ00w2eOh3g1QUvo
m5ekGqXsTy0ppzCQuGKbGaZb7k4jtnPRnc6d3AmVscAblBgDHkqZar5uY9eWXpiGRN44m0/ip8t8
acMkKM9eplVe7dQpaVASXG7qVo4QNBMoYxZxSqmPnMyScWUbebFUdU2e2w5I9v1qnHu57JItRYQc
kFLv25VlpNDMZ1Kp8ajE/VVClfJIU6UsvNm51tRj5miSs+4wF0E+KAkQuf8PXpva322I0WPN+Ye8
GidrT+XrkxpTvTTz3CRs2P+q7SfLYBuQdo+pgF5fnpqVn8A+NH+Jm4fbotjwFTpPx0OllaBa0Tqr
rdAKKMotPD76dcHuX1SC6bClCP5da3k6bCzLo/nBRoqKfPxOILvrJEUW5aWIwvQ7RxQT6T+94NIE
T8pf0WdYVrP3ODik+w/Nf97Ay6kGXlFeinS9TzaFUvL1/1HvEc6oAuaH1yQ5ntaepMzi6lvkZpLY
ecZgqmcZaq/cSmaCKlGZT714+hpNdaxMn7B2Ul61HdJ/ukiDAIkwXhb3GRMFKE3megD+vsGd6uZg
zGqmHkM/XOiIzLowTpntOysRsFKYyZkcFLoZGLOzVBzIYmucvcsTJRrHA9J/xusV8WUqdvM9XJsu
AVyn1Ryi4R4tPMloWtXxL2NHd9AjWhHqvjPDMkL+7Auvn/K89/NL+5EBABC35PQIaPbEEYxSnA+6
uuvcw92d5nY/P/wyAUq0157F+0iacR5nVzzBcaI57r6c8BD477H3qPm6cim1zqQtKxH4KPNVlq0D
kQfkFdltt5KxWFfk6sKvEvb/1bz6eH7YYYWWtAIETUhNg0IBwbqjsbRHixaSlV4jkG2eq5diY2O/
dVvTU7hBqLhOFkqXZPtzN9FB1/zkm2HwKP2YtQdNXAaR+Ar1GCvZRcNZhAPMzYvtFmGpMLo7vCGa
WdOEMx8u0OLjhxueGHOgxJx2bEUPYPAmMB84TtbHCS469tb3Hi0uZ5TJDLXQGTC0BOqrjICvCkb2
TLnu3SNke+FZxdvSWSAAPMPoTCMZr4cc/3vuNvAXWm758GTDlO5eiy2Z9JjXXjyjvptICOH8D4O7
9EmvKTZvaXQ2CF+e2xy6bQ9oZCkOTzi7Kq4nLJGWud23whSTY/ALwGjVKr6taJsaNlIn4a+wOkUx
jc055hUXUp23O6miSqlxpOtSYHl2eeGN+wJErJdGAMFkII5lRjAWis+S/oifGNuyCUDiBsbdURNy
X41B289XD6Y1yw26qOK3BmOuZ2iQv/sHjspjBie05o4WOi6Y9fhRG70VGfLg7bbtlznAlXkQ+T8J
ms95jomBVt+B79vYui9VpzoV+vj9PBVVj0t2w7QClvnLygNJ5oiS0l3S/ARHtPvbf9GFfmStW2zf
Z3gvbdOXSgIhw03rX+8XKqR8hQq5V+PlUyPRQzb8OKeQFBDrxBaLtIhB9mZQUduj8Gx2PmTUj+4k
8SJLGaJCd3EvpqzBj1R5dVVJ01z3oP1TWpQSLsinYT0uJuFwEl2FWRVAnEXnx8xhu0czH12T7P24
SVeB0UByAFXogsscphttydQD3V8RTBncIMruPPFIXjK4UsOvMEQowIckx1khjStIEvm9prkv71M2
cLewcY4yhwDrtmZHasVm092gKWbv3OZu6h4iKWoIGev/gWmwmsd+FoF5iqC6L6+el3lBIhkpOaYw
F/kI0hwN5LIOgMMWoO37aGrsTF9YGWFzI+t3qA1eW2QsenSsN1a/E4fIb5jzi7UN1wTofbCVF5Jk
uV6Xv2YZLq7UGKCz7ugIorPvZG1vxBc4mbDCYtIYFV8armTae9AtOTuyAv2kq+SUTm/3nuzbQXTq
oVbg9MtJcdzv113ROtRgozOuqdP5OxzGCzwxfA9abj44E6YQk0VztlLC017/WeB3egBFXStOHZrC
BqPffqxU5oZRUQkZ8e1jg+tpUH4COKVhYX9JkDxi8nh7XQ3PQzzI52ziPHHjsPic6j2G4+g++Q71
H6YlZaTX8FXAqq1I0J95bovl2fPfUfXNm1YL8wJdFgmbNsOo5Bn66vxGVB34myLdvntqQmT2BNb/
p1zJ/4b4fryOug4G6MmWfNmKCHTbofmkk79I9HnXw/zXGKcHmHiOGESKbgR5Mk4IJ4GlHTwtNo2a
WZ4PvKWZ9zQ/C6JsVizgfU8Sx4hAXpE/SGJJSm0ugJO/QsD7eBeFtmyzzirDcB8EWAsSu01aTd30
0uzknw9Tf8uWbgfUi6dn39al3nlbr4rQv2GndunEIeTfMu6yPYHw9p0CY8E4Ih83dA5wnZy6MSLx
B5Ws2yaCBBh4/Kss6tKw6Prx5GbOGO3KHxOHYiQdGJlcoRlkjMUwI5HhD7254/hgSCbw+XHWKZg6
FxonzboqiMqubL1xuxJSbcyqKhBxlemB7iTKxq1If38XFWxvb6ncDtgRO03AniLUDZlQrvWHRFjh
wJu5HqgebMjY6YLLpe2m6MW7nwfU8m4mpL2Tic/Agge/CivJKtLwIDgVZCpsLlkw5jKXTHNubAZp
3BHG+ZLvn0zaFQQHSRmDQ9VEA1HoWvzWFhJZTNjLkHoWLV2Fy2x81Q3sP+dt8UAUBou6/BDRoqgn
JkVGHy6DdorVT4d/tvNJ5E26VXmSBZbtM9pVIN10OFPfLF0/wee6NTEMgxAYVBnUcfqHeqT0l7kC
ylVQLKqxfkFm7z/UeCx4FQunHORulYPQmf9tQtUW7e+2L/H7Gi7QODMTbKWCv1ymgmJhFaUMIfoR
+81q/wFlWL9q59Lc19uW6KXPrhjiSPJjIkSrEAqKXoq5jdimM/mZReODud3vQiMZ98Wv38o9NW/X
+bERXr2VxJyCl/JWweKDXPTlQ93U1mek+F+G3Boi/Ya1I1bTdfWMxJdh5x/AZV4qbEKOXBI+iw4P
+gAQjJ5O1nRZDZSKR3tYFGGmP2Vp8S+0Zq+nW09QoLDVF5loAtBxM/KjO16hgDTEB5zpQICzz7WY
6MuQkZz7cOtAc35iTGSn0YBl7Q0cCcYzZzWCJRVJy3Cqpgh/oro0ZBXvkY039hKoTyLV6cxfj+fb
nZ0tzyuP7wqYohD1d2MrKU68Z8rhxlXijdSvrtUnVEX+cfdVcZWrF2/GqGeQmN7OoOBVJqQ3FmeA
vIxj2oO/hFmtCRg3OV1JAcM4dFcupPdUZMRQhrKurh41aHIl/K0YwQUdwXGcb27FZGgS4CrtC/se
dlKjpq0EjxH8LfK6uBMz6SwCvg4pP29wTtvEnBfNXdgte/Bba03VCHIsdHXq4xStxPo+OY9tv784
mkM3QsvAEMfMGqwTNkCk+afyVs4wJXQsG2KevIXVFeznFIUeprlC7Lkxk5P6LKwTGvF9GPAth7f8
2V4XMpGvs++qCQpGBIDLWL+ZjU0dFVK9OwPJJufEx7EFE6j6+wDy1QVC41GmusC2KVPyN/DHOQYr
eCp9PRrur3Gujuy3yFNH1azer7se+EMoYXfifEm+bzQzwOA3FuUPOWr3HZ8o535/VX/57Z/QHpuL
Trytd3B33tHrnvZ5deCGVgSpBFUMzmUgTsroact7rOu6W2LMKvw5J9o2sHTrehYerqD7nbHzTeiQ
+rpe12vcAcWzOol2nqEVTNDnq83NpOU+pftv7zOZKhYBmts8oW3y0KFvZrAlkpcQTvISk8glrvRk
H+1PUcLnkSwHS2oLGklrs3d08x8FYFqB6KdV4HKhUOIoqvBINz03dAi2852QRtIYGShuWRzpByq4
p1GgT2M2d0cNyoU61Ekl4/wbXrjcytULMjMR00dRIZSenA2EC2cdFtpv8/y/gE3j/NOfhHDpStzk
py6k2du6qVE62uTh8ehkDGHaBLP86IQ+hjCs5wtAtmCrPoge7eqhW7YYfTtmaabwrNTBF5oirkgV
epqzyzr6ZYTkyOG5aebVr8NLMfJJOFNpWv73mdnHl1L7Jpf1b603cnTQ4mDf3C9QWpENDzP/yyTQ
E1+1yDXcqV4Iyv08cbN1glDzhpN9aYB7ty3a/I5v3VW458+QArzNwJIUINkMY0JR6/tDBNIyakYW
D5V9tf5zeQzizSq3yTFC+7zSCY2P0ayOp15beqfEskb19HJ4/STXt65qOVTi2MMIoN0IUUBS1zhG
RTc+TdCnWe//MenP3URYNSOf1pFlQXppTSwCBH1STvH2hQsGZ9E0V97Jj1n76Kd2K677r0e4qMEX
Hh4Paz7UEScOeaMG6O7j+A5eHGPUxo4tYYa7Y3FhTfPDRmORFYUHm7Yp5KD1BrTYY8UanFkNhDpZ
4BuPEemqieCSb/7VknWHUBgXx/Wi6X+EbD0vgIXPIEFJhxWnl+Ih1VhC0I5JvG29ATiBNf19Ocfr
LvqiV9oT5cm8mRr+8V+NYvNtq99LQgrIbe26Dg92K8SQ3t1pqS3S/MLw92umlARdkYoIOG4oha+E
OjxDlNtoeDikSE+VJ3H5YNtttM5CQYgQk8wWj515L34drpuzk1uaNnj38f/nwQKbbc9tRhsJoGjM
gc1jeimBb/koGHVMXAaxnzrHaA31v/eegZPeWSrWWeEz+R2TgdNOzpQGbP9c5hBZWGYjBhKPi1ce
xM3uaI8HvshXy0FbhTq8mikPOvQBlNN0wDcIYBJGq8db7KWAmyOTaivQv2q3QMMC1gShlQWK4jwu
awk0OszTbJYqhzSPDHu0hS/DlX9XUg/tesZ5FR3Zblw4bgBS00EUDOqYCPaAuEclHAuY2KHMM4G9
i+GP4VnxJkMV4l3adKoL59OXbdWK/JEA8pH6y+gQZRwU/I0I0HZjfB0lX/u6QHsDhs29KqG/9U/9
O7cYaaKPk+XIl572MJakLskLvVNf26vLCr6sZiP1uhf6L3RO/Om/29VzQ9sSK2rSObUtAEcSdftf
tZ9HcDt4xbInGJWk4dvTw2Y8fP0SIm5OmtMJkhM2jMjJZHfq7VHQlV6n1VRgHLW+At4t8CSr2y6f
wFC4ogc6hYAd6PgFDMxhxaWOKwV+TNR4P6tbNnmuCjo9TaObwS7jSr+GYnnEvQdgVqfp6G/em7FK
0Lb54EWaAMq1NRP+F3wXbKdDI+LXB4A+flSVItRCPQEzT0EAtRYfyNAhZcxlpaMDORldcslOcihl
SjI5B+7wjXJCw10iB7ISDJwxrmvRgh/CQ29AdTahKmafWm/sQhCDeaFbC/ZvZ0CIxhzqwUHv212V
yb09Y0G5B+3azOMuaRYCK7dq9wdmAMOIks+MEkbW7BJoJ2amCAD0REbudw+zLIPs8Ienp3sMDQAP
m85tnneQ9bQ4XY8uyliYFyj/Mm5zQU1e8SNOxnVcCekLE1sZXsQHFwOiJDN7PJ4AJn58+cXcgRVV
TPm5pH7UX/5kPb5adhNiNiJu1PHSFH+O6T9uujFjK/qrbG0KRq5BWJEoUIvbSxJqM1KMXxeQCBDR
87ixpLht7XvElMpKu3fHAq7fBvOAWrYeS8R5LAh/NHvDv9KR30BN6ptghS0bpm+yEUluLp/BN6wx
MngpUb4/OWN3zv33cuPjlbeqjGItnU4R4PnG3mATngvVxJ1lwOQw8klZwBgiXMehVlFGv7u+8S8r
JjXoNM5mFVU0TRChKXbmzpC1kkWFhjb8RCQkXcOtkmx/2a8Ivuwps4I7YdbNrM4EFIZ0Yo1BHjzN
asLGGLd6TkZH7hMwEHnghNPo8m4WOcoz7IvFMytHjK4qP6o30KiYrGCXiAjyt2qKAmtqZp6tvYWb
D1XyzlWLh+ekKnS0vQeNtmN2sPDFd60weACGijWIOxzz8cmTgqbfcfqjnopzpC5wUr3QOwppFEHC
cCwQPYDTkHHNgjgwYWvuRkLvB3VIKLt/aJ7hCOOGPn1F/Od5LZrLZAJhjDUHGuOmYcnGJ1wqfiW6
9Mp00N4GEv532J7tpocPRhkGyHKkHyLiaoEV+b932q3b2jMhkrFbU2dX8MV35ZN+CbGDF19iDBOr
+Mr6J5HIaMzuVva5B1XXfhJGz/IyZgDk6ikB1MnBhleTxffo26SoUAvNnNTwz6IjgVebKDwuaKYK
Sv6sjc/NRgyx0cLFMCXKu5JdKFnubn+OLjrLHv4v5468QwEWRypAdR/SWL9X3qzdVCct3m9U+zSG
huSKhwEsx3b/uPN7vYZEdTQ1NhdGOzcQnEzXKTfMNCIJV32gXmduW8rmG37pAg1nTDCSU1ke8RTf
wU+h/nPYkZx0wZBfJhm4HgiluYoG+mbjEP9UkSUJXjCCTu6nKhZkGojDfGcjzw+keKb++ufxylnP
HmRtx1dATmsKkmA4G5RfJ1WV3SOqVBA5XM3D/ecGRRRU0vIxtIImFT5KddJOMMWNo42R0oJD5N0J
Ghk1VcCX92LCwxRIYA/z3L6iONIAg3LouFI5zB7Im2Ytzpv069dIg2kwS9+ahCaSoB9eS9ZuD6d/
w2wSq57ZQNtyeRFsLa4o++r5JshOU85deUeX0oCz/JZJlBXHDBI+oD1/8H2fyFXkxaB/0D3ySKvq
0a3XOhlGqgAjZiC9SuMEaEBPr1oLuaZ7rjemjHRTPl49nIklccbGR1oiC2S5lZXgqF/Ahu21DKDz
sOQSBuw3BG8I1hZutU+zu62H7gmDqEGW+FN77sdYAzChgFwM6dzVV4QvFUDYCkaZSIQRUziO24M1
2D7kBM1KVr+r9dtRORXBopczhBq5xqKotPqpHXhHUuLHgs/7O5mlvns6eFUecr/5VET32KyMbkZ5
HP70QAM4dxaNuJCDiQeTDtZzsRUWtiIlMs0VEG+YjX+9wN0T24t3uReGzgPMq/8Mgp7xFKwu81Dw
oIZtWyLkqW7xx0Q7BdTy2QJOmZSlGW1E7ipCZu3vuAKTF5/VUkNUR4Q8ldmdj2WaaxTc71pmUqUi
rFM5f01GMVrnf9In8iGuR+Wf87jN8osPLxT2Qc9SKOa/n7bpLFfskvdHz+sXI6bf88GjCYZrWO28
s5xA392nHCzMDjFNdTdXs/tu1qUd619vjGSqKz+Aw8YYV0AFgGk6bRdzOEQfoY1ul85eCBo/R/J2
AxlaviZVo014Yu32w9hG2YQpUEaRyMqvrM5R+uY+KIT2wAmukEjH8q/Q9JjNU3gGnOaBSSzcLjZ9
8EJQXMIqCdgLoq2NOxKizP/z3FG+lzWuZnBtljF6om81zDRjpkLBlpLHR4uuodftA35ANAtM2c9X
iToKsnZG1wFDvPpq0+5RVsV/+93XOEqi5YekQ0hdKidUEHoHnPmVG0VJBHp9ejYSPhoPfKrIypTX
bkVHtu9KTaa1M2YnoUa3jI9xxqiUmQBFyCuWLiqRAcpHmseIAdoYkfTWdp/yfa+07fUSPx11dBAf
d3MpEkpWtCOho18sTGG7m6N8AM4Pg7Lknlimu1Mg2hlzZ2E9g4d2d4PeRd4EBVG96W1PuUYLVzwE
J0xcxadrlyfRz74IbVKor1r5FFDCDZwX0Tgd5wz+7/LAeWbEniTZXsFgTbI5E38T0Gi6F0TtoSv0
dx78KFmFyk/DBunwjOsj2wPigSLjbdA8/knJPliqZSlPq6HUIvDu6cgVD+b5UljGM0EhV/0q1VNn
yh07+GfkRkiV97/2x5PcnJarzoHYBkwkHxwzo2v2b65y+IeKYRULlEgrn1atU00cFcumi0nNaKu9
IRsw2Wx5TF9IyGA9pSthjj6EUdH53FS5oIqNhcP4OOHvwSScrnBqd7MECPzkXSjmAerF8qhUP+gb
rakkP509xu93VtEQhJ5s2DuJ4TyrNeEh8gdEPrj9PaBuOEba9cAnEVaqSKzfuVDS0M7gB8oWu3+p
Zrs6xfhOOTfsjwNyQ3uZwt8rjr5aOaZp+QtlbaUHaI/zFmWO4dpSwHcCLiH2wWdvCprUgB4CAHy2
gBPMMS3o8Tb2NPJzam12w2DglIxD8IVGtCmslu6/r+vvHlPr7r4xjF00ubPD/WcBmTk/vYCwGL0P
YdFjHRDoLBKEYBzsd4ww/6LyV88OtL5I+rUBLbU6hVhMHYTaI3WQJuegROpd88mlN/CKPK4zmq+W
Q/qWxRmAYQnuHQX/9vBl8dTDJfajX+M2PiKfGfR//B+Mg4N2CtnJup6UPMFDYKDGPewTbMJorRMT
mN78IN1kU+W3c/2GOV6czZYlJ4dLyyYzSnjwXcPtR4bJdlSA+CAsmCSvrzn8Lv0AX7vma0aDpan0
uzq+mQqhAPRvhR2aD3VpRxgcMqS5Ct4booT07ro7v+HhrWl1MiEWNMITMWw6aNNhxHncaVep1SDF
YUYzzz/BqlVlTPzc7HFIsztEO+1zqDZvE1RgEgLRnLEOj/xMX77LBQkilTfvaVrV0pPQaKkZgPW3
NOi4cjoAcJdeIG7vjkjjTgLR4otsS06YUSn8oVX1hXbW2VgqeqQTeuPF4H53kL5dptPBEt5Mi8S7
EX699KGh3GpZsjt6Df2E7uvJGu81sEN4wqP8dixMhHcczC/BAZYiMFl/5+3ZuaA+a4VhqxKWvebg
OftzV9b1tUmerRfX/30z+HOXQxwZeVLuDvNrsZvJ6JQAwmhyJJGcQeHzVm7bzjBoc55gYCJNjMHQ
kiLjc+1aH1GhiW3KwX3Dz0jCsktumee55tlCCSZOl7xVdjnC1MAWuFk93eQlc7mG3iaG1FJeZ4c2
bAWNL8sebNJb9UNcXESs+Q7DE5+HUfIt3nF/FEjiQZbR5lgX+fzup3+JLgucUNOFaVHpwthKkkfD
TiANlg8cUZc4ZVOSuZKzcH6I6tCIvcqefxfZLBAJWfkmtukE3hEE0LdYORWyRBcH4rtpDeJ4gljA
DWIlBfhuI0D/DPqElSlhFUe86lx2VIq6iywynrvyIokzWOq3f0hFJInWfQVIn8kU638NVv5zfP7L
KMi+wgYqJyZCpRNMU5N57JNKUDiH+bKEk1hyEsdq1nm5YmK/I+Mu8OV2Syrk/6fo7anF+Bc2ytpg
Q/9GuoWYP2RNYKw7nN8QFcWdlqcSdAZEvcQXT/owi37t0vif+/emhxNUSbXOboMp3P+BkTetMNzB
E7kUPmL2Fkw0gRnFUSUduXO9c09RNrizLZ8xqK8SQHQQQIF9I6lMqTKffohx5YKeEmYCjbQuENUR
U7wXbdDP8ksFH+l9X2r6UFjNA8NcnKJxT98B1OBu2VEAjRYJ+1QdJ7BkGwqM59XicI9ErEB5HmPI
PMcCaGuHP8cRJoR36RRmy+TkhwvPJmTsKcOfgYfZPXbHr/uz6qnIvlXglYf2KBebAdfOhmVYJqr2
xJT9Hw7SVUS8HazCjSbNi9BOa5RXbddcGRp5EtTvSBrvo6J0l94egPVOZ62yA5dt5cob9RgXCYac
7/zBNliKLJnqWUcpRayjzHnfb/TGf7wA0lmgiF0+4JRB3wGOHMDG/L9+2dMTsW7aJGkmPK/EomD0
NAbyWAJM9yQWxuHp8N65pvNdT4CD7jJuz3dWRshnaEcpe9Fo2PWntD6woBQMwkCNt3eNLj91LIRJ
gMg/pkH2jflv6721hDmHLAvFPTB2DUd//GYq82e3LTx1sGqBNti1Q6piltjOkjO0SzWhe95ZoeqJ
ACF0MfDI+gPBBmphM1cOegpALtslFw7I/qhsXu6rZAP9DVFlul3VxV5y+DTdL+gsNA/UANMP4bdZ
c9Vylhcpav9Kyc2DcSLzB9rXu0O/DAyyLMPV0UkhUndxM2/F2xZq4iAoeTYraFjWeK5x9ivXwbyS
NOWvnLY1XmpxMNBbm9Hg7l6blZrPlv0blr9nqcz0UO5GG/faPKIQh7v9P+cbEKn+BYSCADwMv6mL
z/BnsU+nDIdeVKAjbptPbBX0oLEFRKI9syJ30P44Buzw20iYQr6L7NVBBV/m7WY7NPcZ/V4jfx9U
YMap55fKGo9JU9Ki0cvuZzNnCZPqD5uEtAXYsEy47KCZVueE95VA34DZU33Hj1UKiqOX+6Tio1bW
7juD8gu7HBfkBMvO94OwgHHkdhdyTDBOBXsnK+7RwPCacp6Uq5UIWfnzOD//apoOUuYn0jgMRzt0
dg79w92/qd2OZlJWmRLvCtzxmmgroUWjNQiFKk/bgWX1CKvZ5a4uT3FWbTAGcZRmJUBMVaV0DMqC
hbUxh7n1oVW6OwrXtI41CKRri4VdwbymGtNwPDZqvF65ljWyCnUO0djKndSV6ZrbJ/Cc2xg6J5Qs
RM3u2zpfuOGw6hR9qvfw7FMnXIa+cxNs7Y2qITZxXduzvWAEaEIdR5H2OneZ0UgOiKJi00Rv83SS
RiDJ21NCyx9RYZ1ouoxr9gSAB6soj5jbz/SfMYc7o6JfZ07t1j3CVwcpqErB8COJVtYnAKwdeZkG
DNjfDATbKNnPmYVsdM3GlbVB/21YePor4gz9BKLff5p9ki0ghU2lIepxiZwoWObgYs6Lam4BcYo4
WEfudDnWrFeF+RKlU7pIwMCSYwWfNCvd+Ph6JAyRSRqUM/yJ4V3E154pnz54WtSGrMcyis4NpAen
EyBH9rKmXi+VzAoLTcdca6Trl3TzCZbm5bxI6DA7Qz6E0nDmqw2RufXep5bzgQQfK+en8WTfYXHd
Qw+dyaI0W1M210aAZcKclzaoWX/XxtkKYfNyb30hh6CZd/f9RaYRDgmJtx/29o0ixMy3hwj1726i
9+cqcPh+gSnl1D70jnVU+b8PrUZqcok5wi6C33HJ38b4QeeWe1nYN82QwVwu1T3VSX8O5V+1OKhe
Yf9I5M233fQ3ys1/XIv1I8XDawiIxdLlyWdanypZSVR02v80o1zUrH1Rk3QXsOkoKKCyK7UiBRiT
BYdc/nFuBv18m66RTgSyi7mYpXaFvayoiNtchHAx7Z4cXgprzmhDI2dK0gG6838WXXg1Gh2JP+eZ
yuy08hBsdjV8VIe/w74BM6G7rY5Xi6eDjTxYe0y3G2hIQR8MZG6ENx7YSdDEUVPcl3elIljP9dY3
giPRZsvZXf6WaRimc6Ew/UAtKWC3QH7CJZA4VVeupnDyEOm28KpS+N3i3RjP103ZE9LUip6bK+Qr
gY9z3Gm8epPxtTFsW4VehZRVgLnkpn+WI70TpMWggfJXNCcXLw4081lZHc7WJJVAXqmbKGpsDlzj
padtcoHMVHduMaJ2Nv2SnWJWCK+kZZ5jV/Xhy7SqkLCZoCCA+fNuvLeKoFhPtebmXQKkS6NWStw0
xcwxBHhWKVMRNDUG08rk7tMe2cBqUBf079dHH/EjZLGLSg7ftxxAgfqw5BYL7zxWJYJYGu3L+3/z
w1Bp9nHdbZ3a1/Xx5iIU3RxfHYDK66uFkzWPnXW9UJbBy9QaUPu+A5jP8XKfu9BGWy1cn9rfAR9O
tDsfTSdCemNx3yVzYPEWcPLXp2ApjGUS/gf31Y1hOX78CPhM4VgtIkLR++Ewbana+9F2ZDU4soWf
qe7TJxIeT8Jeg1sPI+1AUgnErQolXlul1aZDsGngPVUThJTWM86zua5qxaSGkceKiftBkCn6LOdf
LorFqmgDyAKWVxgqb0sviOp9qHejJjQJaFyxeKLx2wLejZr4krCwVX8EUKqCCl3hqdlTFw2g51r8
qfauismLEfBUdrA4YoAnc9uIx49Ijv2zaKdrt6J7NyhNAAqp7RgGl+zpA/X6cp3ECusVih3xHTJc
k6UlO9LroCJBlhbEvfCybocJ+6e1qQawxbxXcW8n0MXWSEcboqkCMmGE6Pt9IU2HhzpDWoDl65Wa
FaLzwwwtr3vi7Kb62s9iVDZf8tP38YM2QhqiZxFABebiNXSt5FTNFFqrzh/Jax+wJvPXp3Dlwmah
XBjRyz0nEYntVoiUKIj54XOc0KoKH2A8ksrdOkR1b6mFxezFPHGwEFldzdIMGTRz62E8wL6UI202
mhtX7zS6mPB2b76vc/RTKjEYrV5PJHtv7LZgocQhr599gNG9TVg5d9/6lIMW5uPsYtDfRY+1mzaZ
N/hTn/89M2tpm0EzHA3uyTdRhpmnsN32xNV1l1mXsgfkBykSCWhPe2Vw0qe6mMMHVUKeYCRxsOWy
x09gT/e+RQIGrnztVMc/fy68WnXtXFEPBHAAC87YVZsf/XYEc1xUtD9wBUlGCrPUbgE9TwAphFtW
c/efr8DNAjN/2KZHHF8QjBuAHcsVbzCtzNlhEEZdnRu0y5Hwq383VqhL6fEMI5AY260t9AdokGBt
OYbdKycnIoBNYg0zjW4aOp+xuqbg8y4yOfSzzFM9oh/xMz+HuFeXoE1S6mUu1zZF2GLGLQT3ybBu
QQzpqOlcp/UO54pPeNx8yNew94abncNgMT22m0eNqTY5Ab2A8Bj1yINCU6UBr+sgNNvZId+xnpOM
3qnOgU8+c2VBqMKf7b4MDBu9Sp6Ox98AVRbX/aiuBGBz+sdoaabYeGcGzGdreDbUGOjmg8O3S/pU
qx4B0g2jkQKf/RTnqwAnMIO6QIcMsRw8JQlega0/Y/NlOybl5dMoWS+6ePgRORWIsI7iSeM/YnPV
oSVwKzv8ryhuodgPvFo90dej57exhtmYrTLWJwc7L0T543IN/1HJ17Km7TjmhYms5De7qFgocdcg
veKU1Ri6CKNvj//ut7KZ42HlEi6xq5Sln2DRlyCWw16zGw9vDsAMdibtilkt0s/6jB1nr5ErOZqa
W9dnuqfHuIx7uA0dRa1vc+nbEcMz9DBg998Emq22hT11bWvQioCpujx2WhlQPRs6/uyHhv3ymKoX
ddFytgzaXGJZI70pIDhOlPwTr8VWjU3ZlGsJvdf/ioRCA76wNlke5nOz02azaVq/KC8WKOftovjs
O9184LvPWCZBfPCkYn0DBN0jzmTiG2fUvq7pADkDuU8J3+L6eqvLLd14qxM50bosJSo/WX6hVgJ2
c85w7+qHk90vMARj/Ui+g1idf0SJHHZ+OHwijDzokRIdq0lEWXU5BBjtxZvenJyZ3X1RSqYCq+/5
prBc7Pk4GKHMjbBVBYcKhQmQVsfPAB1BB502aclYuIsE2c2+lE1VwuSNdWOZV7Cx6DUn3PJT/N2B
dtb99swTUVAXfKwvoVpTe3x3LvXi90YdpKdmXaZzvbLnrEr8oXZXkj2uQJZ1kHun1PG776rp9eFn
zzccxUK0V4EDo4j6DH10++nOJaQbHXPr729c0vHFn7OEb3g95KGjAnoNRaUEiuQqfsJGqPLNqnw/
SjLXAYDZQi4T7Krg2v80YiLcBUEAreW7FHO3IAyvjz341MLdHPqV9pQvzVaiiQQpeHxMWoCbsThm
wwUeGbwW4DQAVfgLdpJ3qA8hOrDcKqDEOH66zzUaOMwaiaNYtF28i2VSsIVkhpIQsYK5GfG+iz+S
R2LFhmaXgFf3LwQrTKrOfkDVy3aUIGbELfUnn/Yam/5kbYYtrnQrlJyi9bPWP58mW6kAdm+OUu7h
s6TT3gVM6oEkApUDP/dUN5ie4g8rGYnd4s+vWNJ4XJk8lnsdSjW9prpynM3szjxYFIvR4JmNHtlb
Xu1NLySJUvi5PxaqK5rEMm/anBGRa7m+HOrH5t7naC/YlPNu23WrPUJAf6HCtoNPxxVH7Du2HKJc
W05Hm5uvcJg4+qC5c4GZk4iG0RP7UuXY04qJtf5Uols3iChqMWRXiNRGGU0FeuorYYTNOsQGnS3v
sL5q69v76rMFx1QSqVb2/6Ncoc2G3aKbrwPix+OguNkQh6zLk2DZE/qFYbTffGUEbDeD6d5qIDNn
aSQJERK3Ekbfxtt8V0GwRz96xv/BADKL7Ie3ESWLubXycABxBZ4lZ9Njq6KLagDBfnmJzynKiK0U
E7V98I6sBb4LYynPoouEX85BlweFu8n594USvqeKIJZNg+yZUGJMYvCyQH0eV+i2O9Tzb2X3eUle
1SpfFvz8QTfYqdaQlSAPKMuYF0tGB5QZH5sPDLfjqlvCUXiEC6jFrgzxfLbk/JZwLa/CVh56nSmH
KEzZDkEYr9vD6Be4XmYUeV16YSCFc4c956eilTnJg1ffWZ1LJoBMF03QNpk/d/ZbhxsEK05NQaP0
8FQwNLe5cRHCE+VdCzo8ybvuEGflzW6WikM+agXDAW2Xb7qq0qh6B2iHXaAy5xWJi5YYPCkZ8jjU
CeUno8ozMx5dm1YbPyxdZI7QtD8babvp7dFAxOe3oxUSuN/p56BnLseF228xVgPRrbgTWnQsXG6Q
2NB1GOpoJXmVWxQ+U3rCmtCmfZ18oCkLtHD2x03CsozhcCzrJ+WoP9HA4J+0ilD+Jde1oziRLLPs
XcaLkHrEI1z+oA04fR1Fklwy0xzp1I29T9+8lJr4v99XuKnCfDRPwYPviBG2sHHZl4Rl6KN2U86V
rw5bi+WOJMIbcDGUtlddXQFqWkAFZkH0KptterVNK88URWo3ejAB3pKEclJzidIQR+Ss9yHcoVQY
uG5G8P2c2xKAKazfRTI/ua2zoPTj1eug37CcYRFDde38hNd6BqDqUuYHIAa1PY5PHPmS3p8+X5/j
PGYRMTdyrSJFaesRCBDxwZ2Yn4xIBqRt1BVFAh9pBx9jTbv8AH+245XvV4UZCJwnQkE9snP65/QS
E7LGvPCT+XvKEz12Kq8dxXBW6XYajO6CeAZDDE7h217ph/Ix5ilWiT9BibvKH9OIAxH9J5IysP4o
1O0xe9Z4xF/Vu/6iDYgipmr1zqDa3f4X9fVAH0xESxtMUUJD6dcTuXbboO7FZPlyVuHolGpmT0Jq
DfzrAg271BEOL64x4/jlAr+1Pc0H4Kwt81AQ4eYIs7emPTt8PPlL30sPxr7g9yGoQ1WuY7FqiUKM
iP9vzwwhtZGEMKOgryD3iQ+BhuoGMjlLARpPpLU0WgOi+uep3/BE/fkaGXwmJ0+zlThfQ/U3b3iZ
Sepehnmej2FPvpgIe/ZDJhj+tC0TXrzrbjCeEML5c75htjkhdLTcecEyKKu2HUh8Cvuoz5z0T9gu
C5tJjHC+OW9vusKaqINoF3dAQqfCsPcIRnrhhUifJ01/a73gAI3hlklFwrxrRvp7aKcxXnZ7/Uut
vC1CBxILyooEqnXCEyCKgQF5D5uG/XpNYPlqnjQWQVfn7yc29WFKQa/Pe/DJ14qcVl2p8fC96/aH
x8kW6aBPppVsarVe1Y+9kmnGlch/bAwZsEYmp8TPdxlSxiZTLUeSEHXum26icfoGQwuqG/kOwfSH
Z9K/40IsKoT9aYlbrSygHx1Qg+aWtZFYPzAKLreD6HipMaKwqoYxGx5NZOZDo8GlfMBNXSoFNWRx
ApvwHd86bJ1p/gK8eFYGhpL27ccAL7LrDWwTF/qotHlxnOwA7qc1aRHNMDnmUegfzlP1fOzFTOPR
IOmx5kAkmgRz1TGjEdau35xqzbj04mTLsKGPJkM0Qw09lFiaaEj5sIaS7gSAuv98oIt70ItsHlun
TjVO+8rxdxZBedu9fb8N5+FDbU2lTny64dvIaRBcxROStLQhkp6pzcSHyfG5EBUIybYYjMH/cC50
caH/F7AEyWNDhVlHVTE61Mebz+l9oqRXuPY5GYuJbSyU7LeRl4AnHNzIEya366GV0PSh2MNfGQic
wXBPZ9j/9vlcvogCItO6GFxVT7z7ciESaCIhN3WpUT6WFcylxrH2URiTj5/B7agTuzInMO+lmyWX
sY/x8cjBkRBXFit58joXTpMmLFzpeWt7+7bp8YvGDONvYUMliy9bQ62apg7SxRRN0ErEuOGGtiRv
vyblk9/1RPXZyE9KDQ0Q08pAfR950w6rDtcGTx7Hq0r75Je8kMEjf6yYMRmzyxZByAOLQAGsorLJ
g5hHXWJ2kZt3k6GM2uNBKGS/l2gkwD69Vw1K09ij0ksJ4V6LHhiKJ87dlxIJzhFFTGHD7MgJc5fX
GqCijISkvYK17HPUFgBjrShf+Mbge9z+sTbte+N6Bd3GGPWLnVIbNXPBdZTxCpmqbRPd8Wg1vyeB
Ex/QpVnHhn6jFlsl0AG9gtGE+00ehtDLq5/xqsOc9ij8k69VTG0qRYIP6XF/TPmN8dZrMSdrhcVP
nzlbWdCAqqi+l0zLBLthWRea0kiY1VRvoZks0OjUOylaj4j1fr3mbUqgHn5jAWhdaE+8CENFBYlW
vOEHnq/j9KNhflwZR1cXwH9HNJ78m45FiGSYk40qB9piow1xWpVfJb1xPI/u3nEA/5DhPbcVxWQ1
RWswEHUacodtytaWaDmEnFaNQPwAPT7pvvhwGePDyjq6Y+PyO78/zvLcX7vTsT1PVo05Ry/16CC0
zMq3XEus+5IovWLXP8kyxIjNjXCqQ2L+CXIGJa3RAiy3ZlpG5i1dDRNqIt9R1U6CMotggVegid6+
992AcAOqxBag/CQTsOkegsEiqFyndWmoK28yTO6WuRqd8Ray9nyOY+B1ULZmJhrXyHAChx4Wveq/
ZlYNC5Vc8mWOQAN7zHMyXy8f5k/dB/l9OhXkS2nioSAW3EnkurE0sIxxU8DDwVS1TFUDnFC1EQGg
KS7GOLDoMgN0GLYXwvjM73jHpD4oHc28LI28DGvijFKZwVx4QRt7+xDoZtGuYlcf2fQLOAaNo7ZR
idQFxwzb44l2S/1qwySZ8o57kauRGagHjsLabklEyq6uJBpb0kwQYeZfxo/y93k7YnJkqQ6WNi8s
yahZ1bFxX31bzS2q5Wpj6/YI0MLF/+Iga3YQA+CcYOSrutAq9e6ItzWeIhlfWDz/RodW/lqVskfp
GvXJ7hQJ1k/du39wSrbF+FTRtr1w1YE8crm2EaoLR0O0mbtkxKiUfDSIPepKKCr40C8NANvKMjpl
Qa/wfiz6o2CLvg7qTYlS+zsdXm/UMh/Y/hbEzeeCnwend8nM3SmvGDHaOJEILuuq374fOHOl+ezd
8LMZCNM+yzYnNycLo737Fekf1sYyRPShUb+MP1vw4FyZwUkk6twY9ndclKEYhfQCzUd4ta2rxDSM
sXncS7zLDeomx8mHEkiU5zqOqW1CjXkM35h1F+Ar3zzlpKWAl0xq2AR4RdqlUgfmE3+y8L0zRWhY
hq/e44S04reXh3d7FcxUguaO/FZB7S4NyZtstRwbN0yjST5doIZUrsGp6ML3Hb1BM3GImdSXMo76
hDMj/Br2XSv+U5UgopofdSXDKh/zHoxJ+bHgMg1fTK5Y7O80yUIGBLxmXl8JeQaWm4cqyAysyai1
bd+iRSO7U9eL/1Oc1dygLgho1tx3yAZK6aKrKnPDYAl4DAvKEsl4L6ieu3LFM4C6G/Rz2xQy6EEL
4p8kXsYTm+by6f1c+UbSUHJ4Y8GynhkyQp7XnbdReVF/10yAZNcHXmxXZrB+MLy10krhQlP2oNjJ
SQ3NZ7UTOL47K6P2iE68o43FYFQu+Dc+BgYJOaN4nTuDsTXBDpAFZEjc3fbMhXef7/HE85C+46kD
xy06E5yjwmVcIyWzwsuj7SRPugFvJF6mZxJfkOtIX0BKEptJO9dhvaXUjOv1ObHGB2qRKPBdKYBU
DeBgO5+mC/4qx7E4cxKYQflgurksml8hUPVyF/Y0X3UCAMka5mqKNMZYuMwegZNBntX2KePF9p7a
spegKin7vAbDXkU51PruUCRtXVKoJoQyG/4YQhkjp8JcHou3tyg1vhE2ImihE46cAdwikqIZgNMm
ghbiDz1IzLJRuScvKRDcl0Z3DIy1XS5oNJyWwvmn+1JC5uyGOPUmi7oY1Rwsx2kDrwpr3NAXK+x4
/UdcOaebxbd2LY4Ay0dVH9OpFDsM6HPk+r6bYTltgi3XH158s3FAzYldm2cwjZbt2L7B/+c9DIKG
mvlnpzDFlPiKYFyvqz2lTi7wOfi39QVLyHErbWYejKn5HE+IKQEgeKRABqpwWx07RIG6m5t3nJnX
k607pq42vW7U3OxuPTnEdA7p/KlDiXol3QhwHGoZ23PS/UjudHwJfk92/nJXAekaWWIY2wAC99WK
sBdBVeHVtGsAvc7M3i6rDzHS0Tfqq2zDIAS9Lw6neei/R4olA+oK1t5NZ+BFZtHZBpIFvN7cOUsx
UEGvQvl9VH0RZk1a+EFe8yK1hpcs4/GOqIIpSKP8JP7zIlQaECKMmpMQBnXsPb/7LXZcKPg0vqqK
ouopk1mRNMX7ZhWH0bCYcfGbLUt2QMWYTMs2Uj57liYe42npgBCD8FDh9tu53jL2f2sITtoiOk6w
vLyM0yGXREYDuOyvlesFXEwCTsQpbA+Aczjl2Da6j+MlXRVGlsOiHnEtwoXfwzETD8IAQzNTY4po
puJOYOeSuulcpieAkhoKKKmMw+hiymhrBqxHTHy2Wh2Nfd6QBN2W9jfPTs8qTQGjY86RqcxaD4dw
Fso5eBVUtI/aZEiHt65KqFVYKSRP/d2eQgHKkDHzMnWXtNztlhh2mT2NufwyN0McgASIl7138GyU
1Esk4JR+4vIuF2h8CnsfJRwcSMQEJ4VqT0xQi7zkxk+86IVhoZK5s/xQZXOcrXFy8SmDV5FE96eO
Zk5g4+8BKBw7Z9fyhtckBbCr9w+pDe9peVolHLZM7d/88u99LwWel/KAOOp6KUQXypT5ugqztHn6
6gwGxCveRaYQp2p9n1X46GAk7MclI4GF0syVhPcO19btMJmqKRftgUrSjf1cANjfrAB8BfExJBBa
BbGx8t1WwPRXgr4vzs1fqGL7nncmOTGRAuV8RALFghub2tOkiRctu9phs6ed93mZps1+nB3F3YsC
N2j8HB2qytheSTGhggt/mUlwHQtRNfnLImJUudohDke4ZD0ZQTixN/6XrCjTVte1P6IYj3vANrqx
7vVpFpuOWHd98KxEpIWK2kVKPylJxPwqELzVdPuoEYxHKWc4h+tYGpW2jt83vNmelG0bDUFkKLmi
pd8QVyREWKlBcYysAhgGumEntzFvgVF7wcVpPJzayg6L5eXBqvtDQsaZWJArl5cMfaLOf4wYwR5g
j/UQ8nZyTSGrHc+4PgTZ5WcQgr1KQBFVZxKwPS2v3k98mmb/jgA3kSKFxFwG8P+r681W0Cs47t+b
yJrNB16TTXHepxx2y5qJTnnnR2CKY5ORzJB9pwbkugT9zQSFKuz8vc8Occ/8lj9UDWHlDpIgVUUo
DW9vxAV6tx6wQQxlXrynFdfK8Z/dz20BX90PBH8K5+XCvZLjrRq2iMN1F7+XTzoQyTjraqhXv/d1
zVEIrLuR79IZQgPVKkvRIJue0W8tTIb72RbsTpeXuuDPKJWT2tfMLHV8UirSLdZfUL7zhbe8Z4cx
rKBDzvVDsykQRbeIIDnf6JDBbN+VTroEcglPwLXwmofK2Rt4Da8hrU3P9lFG4nlno+HcVNCmW+/w
6pcs0Ao9Ykl8g3FGrJckFKH5h61nwcHS9Q9n3a2Lc+yRHeRhHKIARcSUzFqFdP52UO1WvlZvgWVV
62Eerb7p/dBdl9dxv2t+eGi0LEY969HYX9iBFesR00pdTTNdc68TRL3svlaWtPOuu1cUgdmKKeSZ
uV1l2aD+6MDEqchYn4DnG9tohLi8WvwbdYcH5nC0/5h33SUjbclQM45m/vUQRgM+tLsNb4ldofEY
myZXE6TLOoPDzK7yx4O1YkoM0L+MrC6kKbpaVSzM75Z9vgUf+ycJfcaKCxSwbnndahkZF877DIHq
JQyD7QCVGwDDstNJUg7Z30zYS6zL/r46CQIth6Df9T/SzxXRYeG4VBUm15Jo/8pP0dskE/qnsqVC
eySOOwbg+PfeTsOnDDJqf2lus8OU9puUFnWRr2AkPZqZwlrit2trdCdCN/VoDFlfgAI/kHDtwB60
iVm2PgQ+Hi5Di3zOZXax+KGdZUJGeJhpPnXAwsOaMg7TQF6HhLiYgsltl0T1AxQWVWKWG4lL2DHa
V5EQplS0WuNb6yxzf4AeQxh9NG5d+X2nSXAS9mBTOuh+6lsco69rywiij6Z0GQPxI6qFzVy7zI6u
wUfGH3Z2Jy9Z+hzbfz4yqZzAQZzzrPXcYRI1kURFZGfSPk1yNMvIPqGEiKuybS/DYsFAAA/ljHTM
xi1lpLGVeTzJ49l/yx4Hg7koWAF7am3usla2qONDuNMoMVrbBgJTl2A9L5QffXrQ9R/rqLUYRKkY
E/qYjR/Ee0fSWZXx2LKsmOu81E/sbQ3WIEh5EHdENFxkQAs5DWREuxGZ0f+7RXhsvNPsdsSniMSn
1ptW2oInxGlM2KoMlZHmnkesUAAd7Lutnq9EAOSxlEoNMZhYWZIHfzn6ts5BnJICx8vHqfSnpTTP
yGb5nqtSgBij2FCrnqh8c366z4EDvg51vLoo7FVq6LYDOQLMV9n+5SWSZnfa1RGrlWs9CL2jpbP4
RutvbcQGVI2SE4jxlBuVbRL/X71g2GtZxe/4yplZ0vvxik7MAtZZQtEfkumHqO5RVZf51XDuGnpg
8sFb/0/mevYoEGtD1scETso+3jpHuqU02eGb0nBuOBOITW+UblZux/HbXurljk0bjOzYZV1Ya3nn
Tjn0/LwpNKhIMo0ibXjFdEb5QPvpkIeK9WFl3b/E6NPSNVohKCZOzZeLnWJwJfQZfkJKUY4PbrTz
I/ZzYij0xeIDN44S+TAqZMLA40sUVPW6kCDT+XrFH3oWLgs46H6GdWtNgSWJX1OQLokb/NoLhK9R
NY9H1yytnn9raY0fwhnDm+paBTBU5ll77N9Y2gq4P9VqLBN514DO6UKHNmAk6wFS1dEDSkc1K5pe
rB/JjZIfCJKgVtb2nzuAGCYGOtfPq7Oj3E41W6KlwgUFXMVaYYMVGMLUBrAveFR9hx4YpdVWqcZY
FK3vZMsOXFnn8z6kuZMOklm0aX4zSSRZ2JCUAUv2zzvMyEN34AQfgBzwyXJKGAHHO5iXudKlZ9j1
loVPTCzmT7velBDfNnVuJPxkDn1LgbZS6jLcvDONGtSJ5VZ/zZWY3em6eAjlADENdY9pKErGgY92
J7WHaG+QQQ0ZRkjYFMfEtlkKmQ+EjTlfhIOt3tXC6muQV+vClNxLUK/eiD33c7rt+9qAZi+S0Va2
OCEzgd6LkpJhHjo8e7dghQEtBwVqJ2qqoB49WBjygAE9af6biz6FPvfjnKzqHK4R9Dj78j/yYkmM
P0VWlKnsauLfNmH/0/gFHbO6TmOYqysr7PE6DMW2f0CqbuxQPXKLVC89d6Hd8fCO1JxvqDtAXM+M
U1FCLUHloEjJ0AafqPs7kj5a5+f0wB8NkUcKC5OJD+G5I2XjwW5dKO8Yuu75xI4nz9UZr56OnLh0
zBG9fJXkNagACYrL4HnDt17uoSNIEoCnQ1EMm2djEThTpUqykeZr4AqD6cvngN6eua/KCoRhgKRu
7raaBcrf4gucSK3v3g8dsIJDR5LLtrc2yKJFnO+GQPIVcZWSl1yiWppOdD/RX2znP2r1pjjQW3fc
Y87XSCrAcXB04XMr4YX7AgTFIxzhukplxzl4qruoieqZV2BnMeLI6+mHREKnJvJst8yEHWThStdJ
6VWcDpPESyK4PVh/ylG9NTtYXXw4vYjBCTAJOaUKkG8mepCIq+Y7fbFAMQEUAgHhuAtdnxAAU2gx
GAK2O9p4/lVumLMdwgvSjpBrzmcXILqDms5KWPcMgHRGI5REwExznLtXW3Q873wNs6h/7gXv5pz+
2LgPktlcMobnBlXE+t2osTEsGyNCS7jRc0vyiOMa6vV1mL9OVNgvcexcUKE/Tv5m4NH9a+whpLkD
A63J4EqQcK+rTeos12EnWZPPX1lE7gv0nxM+b6IZtS97ag4TdcTmnUMuznrT4mbIpHLa9JDFubD0
63+6rhQppoq82CCZi053maBZm1UAoqGmhl1dcBtT8er1MB4im7dZ7a/uH2zEJJ7BYM7IZqef59i5
guwX94D9/7t44JDCgBXqB5jbEUVHGktvL6cDJQTMSSPBzGnA4UT5uygBL9FjhUR9/IZgmAOgcfSY
sKFfCQfYOLPdZI2OiibkQSJz2E8rG5jnCuvzLOwue8rd0yPBM2KNUJcopG+mdCE8LKuCo27jcINi
7NAx8gvy414J5IgjuKvvsO9I5g0wmiHJivjskCMpc1gpcx/xtAhzpQ7Dcp/zC/CdFbrsvY2h6tIR
aMxrWRlYrLHhUV/rlu2b7a39RcoqiSGvZiCdSzuDMxR8XPaQ/mpwZ9x1BoxLR5c1A35VjsDFby9V
8tqKJ0CCG9VhjpXfJlSaRZQzxKUTFmdLX0y2dC3/9h2KMKkLR1Rsn4EPDafzaQeI2Oo/gtIL7wbd
oz3jne4L33RUKIv3976NpNSNmfopWJn8UITXQ1AqqYXIvlweiWbeG9ngcgueYf/ZfNx3l4cBCLFV
1hB19mkdRxbyYoj0BZs9nRlCf9k0BVFeAgPW26GSn4+hvGapfTvkEP9nDed7zoBhoOgYFMwFF/CQ
BG7KKabwSdSjWItsr2djwlbhDiT2VHpiJaSu8YlRVNb/DcnrwTQn/P6KR2MGJi5IRnfOSwyrdQEU
6NckLmv/fFWC/VSY24KkqgsftctdGa76Y8L+qVnXZj+sCq67LFcNkUCav5PI09wjFM5S3HthetK8
jhTUD1hTon//W26IsIIGD4pDiYY/jAQkO3fEdyg2Fnara7iaynjts8Zhi/wrr8m0skaXWkVIB4sn
oNRx6+LMyIX7ZIZgqlmKapimbkodFO0+aTJBjCAjhX17LlIucNowQtwalj1Um1BzHokLIAvSnkX0
7PzGYucdk3atwGUqSYJ3Bmcewn6BNQ55QXrIOUZomioOf48JFvt9VuGqBWa6zKOMY9oo8iY+24pl
E5HMBxauVaQvFl4KwJM1TSUifaPqj0B0I6NXzhHDK+To77N5hQK6It6gqAI6FCHPw7IzhTCTTPWt
OL2QSg9wvxkUXMQ2qHCxOQmqbcL3G7tiWg+Vg4KU9uanL6N2PXbQ7tIWAK5U3wopf4kRysZ8OkOR
RgEVs1GjPve1ExB0d6H5C+1JOK6oLHxVgTmXAgrvDmqWHOtfxBDAG7pPWO+qDv8osjPEqNx3Y2Sm
O7nb0idoYWBCg4hCf1MrH64uR+9vIaALeP18ZBEQGwSnxanga0d3gyJyQLMRtwkXRUgmee4gdEsr
vVABD147q3g1Wq+x/aEEkMrR6ocaTcCTYUBFwDe3MNlxk9PwVqoLSlvZUgqzGpyNyupZTaSQ3usE
f5iItn33IElOVNii/JczOSo58F4QTi+2ZR3RlIaFv0522zgsdBwgWftWwmDbsDLDnipUeBo76DMA
ZoiAM6a5gXtHMFrfbGDVB8zpIgSuSl+TwQYoF3s7hvhSCAMp96DcXO6JSqr49KYck8s+vIdXunzt
7ZashawTSXQcoRw0oOjzTe2b+oWkUWHMXn8BCAl8sc111tWBygwvvZJmIWGGq4BG+Js3heBhkU0w
GVo+H0SjldRKukhqyT91sjltHWWPcFB9eL3Baa0rgGcdhxZurlCHIYKRm1PI2zfUmt92DU8hl/d9
OtIeKw9vn3TXxN3BY8EOMNWCddRSHiS4ceaI9XssgTPAwNaGYznbk7AXHjAqI9qFTV2LMzcfI3fM
Q5/q+HpIemkA3iVQPDVqWjYOBmXSf7Z46PE1R7xpy8So1144KfLh8TZI+dEdFxVTP4Pd0LxLMCeF
V1Lnhu3twp+W2jQ4/91yJ2Pql4wZFVxvH0/5h6dECshZALk/1NW0TBabJ8QQLdibPn+TVCE2prDd
aToNZjhCXmRcvVR00vUGp3t4TWGWnlcbdmQHtkgi1Z8v1BsYwNKV2xm/sLH2CunYVNBk5lR7ytHK
IgzXMwZykS8RHTSDpXITHA9xImXyZcvHAJJ5CoeEAjM3s0KxabsPt7+gExDZBmsBD8Iwwal/yV3L
DITZwY2bzAKHemhF+FXUraX/Xz1bNpr97uQqKGCBv0IpnL05NnDSvLC4fi+rKlyg1AsZR2PR57rK
hK02vcQ0grwZKzp+PShIhreMSBrM9lAgULpO4W4qWyNiAOYh1VBQdeTkO5nmNxwKC+O7Q5uY7KtV
TUUkjZ9oXwg7wqdMSE+KQ/vwcerudOlgnvzTNxh2xiuQKrbSFGXRIf3oMnJ/jdxoK9HTJ4UUbr/M
YC/TjD+3IOs1Roqk70sT4X16hsbDfIAKZuGhWBDmeRznWhmWXNnLHDcPucQ+0BURjIglm1rPZ8X+
RNaTDJ1tUDZuIhK6ZmK7GPgQKef+chqDF9e696wgV9jLAiXTUwu/gJZ2FtCViTb7K+Ow9jXTbSNI
I6e21o/nMpJfJoz2ad5Icwean/zI21hPlzIAKHPUtqWhXhQV0ucCJJ9TefU2tFa6+ISHP7qgqhfA
W+pvEkusJ7F5Lr05rYIU6jhGmwJ2Zh3kgAInuOnarGyHUwRuZUhMLkXmLrYR5Q/Bm+nBFQOZ2Gz6
1nqLL00Iw/8oftzoxbwI8vPKiWeNy9Z5hdzEwLAjQ4OZQF+b+nZUzpisWCfhFJHyV5hhQ5PgYt8e
qbbVqmrDWO21f6oWzYlvury2mfG+qzg6xEk194Yv6CFMCSHq0WNccPx1ttu3ihNWLs/6WFmL2kbW
X48GHuS0HdMWwEATes6aAsngAzEqNIpg0cKcAlUnlwRmZiAaw5KfehE1anuPxY5/KTty8LKdh3Rf
r3ssi1WdeMAPlIfGaGKilpqtvzK22lWZMHIBaKz9+AeVUexpisMZQyoX2x5RqrivwRScmVZ4dHD+
cAmTKUPtaL48DA8OzRfB5EO6wEIHf2eOJluac0gSoAmPIR3SzfHMRulAic1O4Io2TPjvblJnHc9U
2ZVXIPf4+p/3fbkDsZLxscVw+JrJms4pilx5iq0jGUWAT1XgnetJxU/CV7ACm51hiCgQASUCmahn
l8e/m2g4M8C+/9rPFtiLy7SGXbf6K/8qivJ0lH4psxCuSR8oajDCNHy63K2OaSTXrg/jWrCnQJoQ
B34aJ9pydiYsbxuL+oF05m/Fwvmv24+XwWLFPy7iZ+fYcTOefv7gp4avnZTKgt0yiWf6eQXs+mQB
cseFvf/YIuIQjo2pVd6uiWrGxiwj9Pz0jdj7b8jX1vhUXv1aLYoDdO89R5NsnrU9opT/uqpCCHSi
P4gQKEJS6rL5XgAQy9bvIrzFBkiKkqHa5IBSNLTvISiTm8aFk3f+CR+O5h7/6APxyS1RQtOCr5KQ
J9NuUXsfaahoW3lBgEjyKblMjkkr66sX1I9K6DwgS/vpMf2KnWtrEBVc7MAMhySoMLqnmAqQ3X4Q
hCwsMZHfFHyXqNQvtFyGBqUFYfb6AIST89vt1pGC4310zgguvhPQJ4EbN+l1U14yLfBafa3geskV
hT3OKSL/lj3PjD52RWZVWTp5nZ57pGXABklL8i5G8IZBdecq5KCY2axz8Yiv6AGN5TFh55FAJ8FJ
Km4ZkTGHAK+eea0ZNUUHdtAYb/BQE+vwwOQxZKO6KbqxnuSQg/Sxdk69GvPz5CIyrL66tqGuyIJc
QGLf1TEEShX4+j3Op25b4C+DpZzHsmzfCoYgRfklNX9PsTMREf21mB0XzNYPp9mSoJzYwA4MHYW/
hZdDeqmMa18GXmxjGYzFbQuVK9dMP9pwOcldx5ePkTuqGqa9qjjvSCmVJ7Y0C0aL6WKcmPRgwn0a
My6KlfjpD+/mx9dFqumtixJ4/tBQDYjeLjuqqqQRR2z+e6SdrLJDS0xzYe0qmK7fje+W5RUex8jG
Ozr3u2PzpTiUCx40UyjW22T/dGFfT5PQ8lBsMuZrTFgf2MsiR9hhngJul2oDOI2MAcJ/AIfVW1ze
39LGa07yggzwKjutZldCZUjW45nmU6PQvb5Cqx8DFLFdECgn0a1oGYX2PADJtkQVAWrR5yXDGQVc
zHMOFOWZQsE6/4+TYjLEa1pGscPlXN1MxfbweBKfXJA7VIDFyIg5pKEWNJsMZpFp5G6b0Z0C33+1
YhHWwN8h5ytodwbH6153iLeIh6ziRgYoDgziSMyx6AtjTzQosGgTGNb0NYfl2x0cnTsJZJQe8HCK
6X33F+0RYw6jHo1cGk59y8kCo7YJ/ldsmjMUFKr5crT+Yh1DOeVtezZphTOh3+YPn6OMqmBnf69C
vYTNAU9SSqug23RCd4xlrz5qIrgieeZ5R6KfoYDDxax3JP6JWTdcujSe5575V5sF8R6VIcAIjx9g
7HyoO96ohm92RyCx+xlAhvAKq9Xuqxgn7C5/BGPjpmsBvYBhCQBbQNOVzGY+P7dtJ2JAxLaV4Ik8
HHt8yKs9Xn11pjlHbI9ePDmEq1dlbfLOc1je3z1L7Ddj9E+o6rk4OytB3LB4jA9Bp41dl4kA5de2
wUhulyjeDY0I30O2a/KNcs1nOmkJDo/eh+VdKKHLOFYxPslsgNGDt1xAq215FAi9qcY1GDKMBVN0
owQwAV8V9yg2QfMi3skSiPelnPyjqtbg1T2npVOtpW3If++oMIPro32HQuiOtSeDoLVhA1WmX/yW
y7HZupwWz6oi6FeOdlBtCsijCnNh2GempfuWKXQdWOraqS+mGfXOtt3oj/UFHC2Wpj9KPcnlJhOf
WIo2E9EHcy7i/no9esq6ZiUREsmTdk7Er035Ozc5NYKtjZdvDeAMFEh2JJxP7p0wT1GM+CblwJVq
5zVbvmOFGniMYOdGSLxDO4+sj9Z3kQJrzIvPmgGUA2bo6juNkk6bLx+XN07xzPB9Ag3AVHQcymIY
poqMxFMekdy6z9ZVrIZj6v/3pzMZ/AGsOeZg6SoiVGV0E8qTNYFf/agEGjlM6z4KZeOANMKvJ/9Y
m73Prko73wWNWnLUBPSSmTKfgcEmLw3q89AOd9P1UysZuv+IT9BE0TJCNmnLkBC0EIJQNLEi4VRt
KrZyR/nE/vWpW2FMD6098ksb2cnEvKqKALg06hLke5ZTiRBcPCXXWf31XnCEa6AU1t0KBvBpM/+A
+T1fnjEke/5G0sEhFSEqDJCIBqX9ySD40mLs3cMcAIkwdcTzhky5j0vLzqvGVdCTi8S7IgymbjKp
TNQMLYQTkLoNJCV0MwI2baFKASNhb77pTN7Kr/xX+7RlV8JiC5WfCmJFYx7Bu+IoSfpMsFGrFOtI
WfRAJc3qPxOW0iGpCeNLF8UsLu6o8tOVA7LejIIrsMbp7K51el/8ntHztHFaitGou0n0Lf9kmfqR
q9AtfF3SIFz3u5QG6h0MCk2EO+babav4r1/iySqc2r+mFP/emOIJfzbtp/A1bivqQwB+EmoR//2O
cJvy2wiFT7e1TYZ7lnw75UIHPnBO3t5c4YqAnBbhNs5vLiUbSkmzXitha0Uv+IsvIXLQBhqcTw1o
Rc63fYhN1TBxCQtR8pdsOxd5CAtON3Gmrz50bi5skeVi1tSKgoFZHgv4DzfeK2lVYNOAG2Oh1xXF
4eBHkPIUA/0Q8t4dwkphkdL6WlHX4GaVOeL8FrqKLa1Mm8227M39oZCuFp/W+PfKV9Ay2OTDR4N9
mRsGqUZ81Q4SFKWLHCqZ31IwGO1TeZ//PH5VQ155y9gfgii7sNQ1JaJ4cAKxeQyEdLk0GnmOO1N0
IRIAWO+ipcC0PGirf79DYtoY+oqsnXHRHdqxmL+CFs9bMA8V/ZEFr6lw/ZAo+MgKRBhtDEEDM00r
AoXdgI3rES/S+CAqvhncjQnK+by0bxKEpmQ/igqST0hYqp+k9owDScSi6j5Tub2hdCqrVUNYKXKv
3mBqVnJppuX61fOLBlceD158UMQHsZcqHFFTe0pVekFzk/xFPg0T760lqfQxu9M+LwGco3Tb325j
UmtaJB14jiRe3jcwwkEIKeyOTPwNLqRLB99+/wntZw7bUhqDCzyZ1L7/zu7pAJ9hj6BnPbNuWJ9P
+7xpYODNBLMM3G74thzLzHO7KuO+ryS+7v3+AqE1Sf5kyd2J/sc84SiDRlIobodEREkZ4+ED9jIU
JJZ5GHyYjodL7lkVYFOpsNVUGDSkHnQrziwnjKqyRcdkEf/wM7OtvzQH5CVZx37BtmDPHLUh9s7O
RNsDSBSyThV7AHg0hvY13hARxYQJlWDMRV6E2KzQA3awy6XayH8DzKDGU/LOsUmNsLy/IGIg56uZ
ibwf9Dz8c8rqidsR1d6vKtCIyv3xszq0LAcdMJEf9I5BDi7SFxAbFtih1K6Vvkr0t87qYytV06ik
RZlkRuBuXBM4W/L86+xw0lnz4RT7cA/Qh+X9dXiTbf3lqSXnNI+9Mn42AEEJ0aUB3wTSrXlZbsgY
EZ547Cx87XQVff5ChrWOiCTv5+tUivpfC9ot1fPliR+Thi/ZH+mwSRYnlrE700gaoKMzno+1z9IF
La+p3JEVznz/bM/FGfE7DF2bO8EcExaS/FqJY6NBa52AvDmSdy7lRAsZjSeZjNLcP9LX4K2JpfYT
oEU0M1u2lBHicl1UmM9zLphYYnFI1f+WCOn/quJBpQZJ8aCUL9+GHoCCf6C8BfwkWW0p0XzlTp69
g/bdF79rzEel64sVYavzrL19jVH6Qn3jbVqPP42EQqmrT1Ox+2vIp43SpdWAK41puTOVaXl9rM48
sQrbrbxfZlY6/2zc4N2q1oIeRwdACm8Df1ebStiQd9TLcGtJTtNTpOLHtmjRSz90W41WZtoxH7eP
eDqjAxJZlIN2rgDIJi51jQHvK9/lQpW+/r5Ackm3DhWKLXB9vecZe4XTJOwegq/PAVp/CD4DDaTC
1pirF1UjvIvJWZF7ihbQUnZEBHk/2NVpSt2LgLFp/rRcne+hB7U8NQ/mWWQ2Q/uwvGZkhBLbNc2y
d7pm/KgWcSzDDUev3DtRw0j4JcXBXTvSFvS/ziaVzcesfeW/UFZmVOdWY5GFSZ+BQjqi0yCwB7Vc
xS9D0IfqO33XaPmOBHGSN7PEc0wxfXAgbD4VPVmxmU++9mcmslmJG0xFToo34KtwigB6T+DUbFSi
L9GNmTERP/cAUVs8JKrpErAiJT7TZ1hljQ/cKREz47+OKm6cthAioy0I2ZTSVaprfZebnnde+kAO
5qgj/AqgjEOztjQ+2VyHtu2fJTVaHMy4dJ3RGfPITfuQxRMcCbf3l5DTxGGLeH1w8KIMreWLEtKi
M7MGSHaSj8or/Ysl4k8BQFK9JkX5D4CjgMNceV/HZvZdunCuu4znfQ3DUMQr6mjNWNc6TVnzKxdg
gHoGY6cE1l69qpJBBSq3DU+lyEJac6qrMXHTlhasm5eCk81P93wXFXgtedSysshADMgi21v31eZo
V6tYQsMqL3x2T+wlgJ2qyFA/UMyLvw/cLFu0atyt1n8KvA95HMeC5LzyD+eDNpJpsGqZMybwasii
HEvj7wO+fXkb5FkRfZnEEFAKXEKfLGA5EUU1wSIk9IK5RuVAxfDtgoPzC1UKTV8/CzKRy3PfXy22
off6O3imUGMXAN78gwUjrnvJ+K8wE/Mj0JKLkVYdCbjqvF1SQ03dEPRJswJ1H7dQHZGUCUjaedJd
e7bquSqD+H0tzxVzil73kH/F4g69r/bEQlLwPI1TBFBpCMa10DG9i07pP5P9I3a3sfItT+hNzGLb
UH/H3JMIX2TROf2hNBnxXeR3tT85YFW6ySsEvOfEHE+/LqlqutAvNZezxNuuT/8Otpg9R2ck/6zS
LZRMuNzC0cZ+VvC1ppQ7He+3IotRVFaDcaC/+UvF+bDLFomndxaJV8icnZH1Up2fQUirEvBN6RFY
1vR7AVORIFS9ALyFGILa4Dnt2hnAB++YgACMEWPGKh+47tFFM6REspkjQ52NBfB8kzemjknk7pJ1
o1BJJtL7QKEq2ywfOgWP+ia89TIL8Aq7FySVUkQGCZ1Rqk5hb/y0IF023GoD7UJMr9Du8KMR53fG
TDw7YN1jfMjNMtJVHozFVsokUZB7DOJ34q9cpcoViJ3CB8go0Q9cHFuTjCdpImqb8yx6UMOZAvc7
PgKteqLCbG7H+e3fN0EAMmuhfHVUZfKcNc1poRFwF78Lxwh3giWTh5FyikwBVi+g2AD/a4wl1V+r
rZFhQM6aPZhSUgQIWUqdiL8fhFISC6V5+PDHx05iaSNoEBCf6gxgYvsTgcCjLeGhLK6EGAjE4KYT
hDufjJkzo+PXVFz99YvNLt6+IHHxFMyrtMANB5NnOgiXCuOZfxM8WPxX/O2gk8GbpxmHedCTFxo8
ePVJ+TdQfZYB5Z808nJaf6Gs9PApGAqh7XpAhqAzamR9gzF4BqG5eRzUeEmdjgHs4Yq2s570ee5b
ic83RZtaEIJggQ+FbXX2w+OBI/1MwYpYFj7m8Z7i/BitGO9M1j/7OLpAfQ7VN6GGYs/z8A9FqiO6
+BGGaKq/osqYBkdxO6Nt6WLGefYatD0UtD4Vlein6FPJ/k51VgCBGezB8q2m4qZFq/FngivcBiOv
96gaF8lE+NlgPRlLSEr8z5Uc/shky9Z7ZSLxM7EcA2BSqqhI5lluic1RSgT3W4Yj6iY6PqtDrdci
i8lqfBoXl4nljHNyMLkU7+2CmXlCwtSW924WUiYVt9t8fxbEV6LwtfrY1dJT8I1VZnaSJELJ04C4
KRU0Fyf5ybfn7YCf8PopzewhBvISG02V63JPNTzVtkTO47hxIMaimY/+IrxXEnU5ZAA4jlCvZxR7
gR0xCdwuWq/71g0uYZitE2gbsUjnLwzNz7JH0FirK+n3LdMg1abUrXPEF0y6bK/YX074xjEuqQ21
GtwzjXrNDMd6/dx4jMY2Iy0so0QVDPvR+1BmlRVCNt9SJMSMHfq0qvF+ktZ96rW8FWGCiLxOe5/v
Dn4c3zcIXHNHofP3DX420E0JcMkpuATzknLf6cwqfBLkyDZVAMKnzLCDaLupwZ6yd2SaKao56hNC
vu8ohiVbCJnJhsI/6wycDtRfzL1yomPJJ+yHxVL+BbPF3N2fKb35xg9AC73tTFRSx3inGV7Rp2nS
HieONqlb05U4Qu2qDt3oAnPHnd3Q/9VPXpMne8k0D70OVhZhpJbV7+/ltdCJzmP8QEDo6TP2H6iQ
nvtINQBzI1ZWtjJSvug1LZdqPwZCfxLBkAYQPZxdUPk78IujbXw4Ehh+S1qlB1mL1WhNH1hAPKJW
3JNZegXSUQzTVMNoHI6alAvnFguGCiJ6JxGnaDiLKw7+VxePQU97ZIEj41kD7tb+GkmFVZ5SmH95
VYAKD5o6PNqZRm3dRTJPGfaJxtRkk+r9mgcGh3LVoUG/BS3odgBZrqfiKlMJNv//f5TZkxqyS2o3
8z3DgS6ppNFdxJj/9bjyaZR0zT75LSYaM8/IFcY7kEgSfr4W7zx0vaAzeEQ78ZSUqONAY7CZ/AuJ
fyph3xKwGiSyhLv0mfMN59v1AGh/6/Au8R0D8QxxF7U0+F7IIQQjLzHlSHasJ784oQiVxmqIiV33
jqAOt83m/dISi4/Fx9W7xATeBa0NYJVPPPBSs7lQjsbEcESdq08QYHKzgowx56xaJfKjuT3MqQva
MUhu7T1Z3N/LttXiCfSkjhqpb2vvV1KbOBJsKO4RlABJf3iZijtxx76gfTmBswbj6wBndLC8d+fF
gyVSpPjsN48vx5DbE4IA4Nbu+hgi1odiNlxd88Tu9MzXXy0sB8lxgxAU1HZ/8/0L1hUd2H64FBC0
JULPFGTlDlp9jQ9NgSCIS6SyHJQ9foJAJkO9kFdmp7XwvolDePmW22uQFaRXOft7UqgjJxCfzgXu
4fjqsZBuHOPf6/dyT1pqlxoVua9WM5+WJmFoiDwdLkNrG05fVI/aozmzRftxtpz1nkMdJR3wM2t9
yvWxqzLcgql7nLGuYHtXXIUcKBJZydm21fFEZJbo3mnonHvEBGI5g3LjlIYHKUsU45irsoPhW9V+
9RrNqp+iPC5e5fvCgnxRmKbBuUTuiByNIpj8XlZgPQKTe326aU/UW6XuE+MX6QArTGmsuCeiHhKr
zdLSMYy6/JSnmc+OLwZkWN+39pplbLuXDwb4YIySp3oprBta85HSlkyMdGm0A9OtMSJFcZW5odUU
sdFm+n3/Dno31AAhVaKu374+qiCWKnuQiaCAZqk8iPx4P+lU6kpwjFPwrxjtJP38CJiyN1uivp1V
PrJo0+go3yhz2l8OabeRqmivyBx73Mgsx4xBC/y/pYUxXpiLAAM7FUamxakh8wVhi3cDsl0wJhFa
34+7mhCKlS3rmyQgWHVhqcgevAxjOzSCgeKjl/FSAH10fsPb57ml4/zPkMaioFE/EIegRP46OCp/
TPpFAFB8UeU4qmmsVb2YePQhrnxKZGwnhjMgavZcEapommngKCQcU0jhWALKxl7NcwiR/EwYa9kj
gN1C39RNHR0sJnThH0UqmXxwvVJT3Pei2VnmUHnP/gABHuVHZfjiGJwDzntR7FiQCI8DD2CeJEFD
OHZqKdSNzVQ9qdZa7Bi9lioUPB4RHSsGhD+T/Pxl+CiXz58jIeHnu/uMtn601ytr58rJVQ6qNpV7
Ny9VE/58nTJMROR0pHyYpQJtW7JdedD9e8jNOAg0IaVDB6JEmKFZLpWWpH0Q9cunVniC2zu4rd/C
3N//ODIe2XDFP7m1La3a4sbArinBIj5l37UxrojyZ8RWmuoYPZyFv1lu5MnjhpNWoqKafpoKBRpB
zP1TvLCABrPKct3ZQdR/RwWA13u/NgUIwnaPfgUuVwtY+IL9WhedVtsna4WFFoHjaTbtPNPehWay
B0zvAds6pFTHku99AilLT0aDcMg/D6wThZVJxAn7wQoQLGN9ldoNLYReqkgLHsF9Ai9r5kWiGheE
dvtkIFOfRAJWZEBKHOlorZVZOAfwjL0pFBYEBzpV66G7pIr8+CAlYGZtaOrpiiTHEcbaAZQn7eGd
ikiqvorJbn6dWOSCS4JGyZY9ngSFT97ZkRAo7fWUbPSkwyblCmMzT7jPNkH3P9ZAzo2jR26RTl+e
EpNqK4XEEmvxrHfckSSgUfukdgIgwQnUbYaZajnyByydClcXcZL6FexUlwdWBOvbZfAWrNZmfTNa
mMel11L31/BK/IV2qWCs/OVM60YPslJFSvnUp0txyIE6f0Cdl2FGTrmuKjh0uQ2sjcGJX4qEO6HG
QNvQE5iQKdw+l6OpJ3OES73Kg29QhqD8eeOCgGcTTseHlvVYhc5CTYRu+f5GdU0f9yH0DKUcK/20
XZk/e3WcRxe+wRkmh+fNpPbc4Aae9vtsAxTRorAd8zqS2srCEjoegvdxp8qOtWErepyYuybiO6d3
7+Q/3Y3Bj+vNNGIQIP6aXgsXpnkcykGkjpb+O0Ym8FtkyOw5GqVoN22TGX3lNkrrcWiO+i3AQqPb
DEWFuEE4Ux3Q1Rbt4BKnNm//Zs4gkflqF7xy8DeDYHaDfer9ZErRDCRMTuHGKFHXkIXg7IuJgviT
be9Wqn8OYI9N8hoQ7adGbm57myXF+e9pXBAr4KaXZ7IsupekjYo096HZOzwRCACbbXwm3qZqy/eS
/JYwxlOhLQ3weB+IEsWwoH7KhMte/IUEQsr5SSwCi4KA2oCAZollIWBsgHWZJrZqDnSlZO1LSL56
XPipgAS4HGfPqS7VdpfU8HeCS57PsoQI5PwfDtRod/5O5CX0gz3e9iqcue+pT/NnxwO3FTsYCXd4
6NW6M7pf6hqCu1BnqRPFyZCdtfgJ4ncmQ7ZF8T+sQrpGGnTTvfkTVbDDBlzPz+vtXefqXiB9JVda
TkuPABqn910BJbuQGBr1zfvFL7zrs4g78XFxrrs692nyfN8B5idrhVQBnmD6mvTfWrbTz6BYEJyr
Qnn9Xs5SjmHD7xVGndE5TABuBNpkQb70lv/fA71inUH187/pAn5dFYBaWaAzXDo+0sP0mgquap83
Mg/DISYX4JfN6rY2xI1boyMh+rN6iwBWr6S5BXA+JDGUZYw7Kxtgl1kK7yP9G+hfBc9QmJ8lhBCR
yOk9nwQDdVfJVxU1u7Xuvh7CEJ/isDLgpnVFHPxVLlJ1jo1SUnpKCNNDg71b42zBg8TDFTeGUTaA
Kx45xtfytcXoX0O1Oth8a3R9Z2Jc7LIIgMGZx3279JhB+g4wzYqlBsbPemQqMDqPBpDyKapTZZts
J/WtAmB0a4dvJzkz2wmxYaCs0fXM0FwoiP7WZeZB6e9baQ5uMLl0wTN93zn3n+AkFFeGtIU4wUWm
oDyohffbhjaAUSfNKxbbsK16GNDQBdMSf6He81pg1QHltlLMbXRp8ns8Ci63NK6ahUfOIdIGPCwi
f01fEdNVjvWlWVkF6LXJccLsRbuIzZptUgcyuA0/5eJ0612ZM2cKMtVlSlXyYMhSLs8DB+H62AAW
XviT7NE5pdXNatWzWqWH8SK4cK/D96k4wVawfiDnDDnZ2pFnQ7Yn/Smvz1XgEIU1OTrKn3T5CS/d
WYFKFGNVde5fIvMV/U9LnXw2GwZDeAtEsHLMYaWfgauKxCC7QcAsEkApzyuyMmkWO93I/rOQWEbS
rHo8ThnT6/AMAGNHORuPsPVmrA6pLALucd4qiaNWX52gfNxs6rtTzssX4C30SF93ywhhY+gTQbC7
LLeQ0Dl3eB/ndFCOL69oouCZ1nn5SPrjaByJfj8+hFMh3ZwTtaf47BKGuhBL2udrFJ90Wh10gt8p
ChATo/whBmZhXvOAwHYtrr7XqhoDnIS39Y2NRTopDq73YzWX6lNXQhNK8kdBU/zgolWsurMIKEcg
vGcMqh3TCMaxHW5tQ7ObQuQZfEaqcMpEFi3FSqLQNnlRnDEMdsDO75A9qk3oqe7xXcV+2ubb2EsI
qXOaZiJnjS0YMpMHX+WK29mEuBvmFBvE6k59g5B0Bd8la8VijUXIojwyuGUEvu9JkDj+otCdnCcw
wSgvEgjiYEQGSPx34NTV23hlw7HIN78o/9mxSa3xVAzE/HLOi6JhCU4oVyxTn5e4hdqUH/1BxObD
YZgbD3zL0EhZKUcgUJxg1Fczd3tKCyYFY3+MSVzqxHPKqFFSbAzcM6nvcwXbKeyOGq5Cg8gj4qH8
+KTz8NV02M4HCCZ/a6e906vjKqXeQJDxuEut5XgkFgNVm9eWw1u7Ae6kYx5X19d1kgdUOWNvbN7+
MfRElNiHFCXTZvzyCtO7cP6TNHPrcotW+axfYTfXHtCy7ZBqWIfxIxBYsbDZ6lY8G9J1/psVpfoa
Dd0KPN9Ge6s13u/R3FIVPFvIeTRkYL4GhozrzoPk2L1WVQJDsdri9TZ83L/jDpSXoSL1sdKImSkC
Sbgczae+I225iofgZxnYX2nHvzjDE7BknxCDP22VS8/+X5s30HQVIWJMZPJvLjZyD/rg3rNPWz6E
22DhNTobA1kFboJM9Giwn1m/NU2njlHBm0allAEtf56Py88ttwm2KkdT+X3Mpc6PbJDpEPPZeKER
xwIt8BnVA0iF4sVlToWSz+jRUCj8EhfRthexl02VuzrFawpRsuadUo6bJ4IH0QR5xQk68Pc4Myw2
H9kH+7H0Q2NhbiYqF9jjoet4USR10hS6InoRyjFtlrowUAENa70RSKIk5eetM+K5qFogllgi3J/v
FrX7ynoO9Yic1f5AVLwUidH0PnOMWXVf0Qt0F6kdyOUKPsWFL+PyyQmVub+IRcaqTt7ZcbicDfJd
dENNyNpz7xwpjaMWP7dGNpOapyOITPaJaIAeM9INzJZ606C0da/nEsyAGFTu+VFqLDu9nsKiEOXM
OsFdBG1cTSfh/C+SF8+Btbqdd+7RtdpzpsP1DwgjjLICPcxFx4ei+1solWtmNldMOqUOsYuVFG4s
8bjZrxplCDd6l0wR5hzzk0Z3tbPnFPXib9B4aQSgKs2C0qXaaMf+A3Y+XweiBxeFbX1vtLC1ShaJ
8bmIcAs/ynaPlxKTUEo4JICEJMBPH1pn/sTGGx3bir2oFZQM1zBiKBwq1hW0YNo+K+PCpjwDD4m/
juKZJJcrcXQTUBVUeSjPyru80WCMg/wfLW5QwEPDrS3TvWRKep5sPHg7dkWqU5E1pJ+sUio3Gd5k
hbASeRQK7tFojp3I4lXN8L63Pa/F2cFu8rKi2JPYfzaJW2t7TZM1r5ma8BDTDbZGAwYEQzCUor9D
WXz9wn0dTVwwWcCdmUps74Hj7SLQelLb/xZ/OGBaggVplUDxUFEQKSApeOjErAmetmj02o35SGIo
kf7i2qM8b5JoHXCR4E552s1qbEgvzODn1SKdoTj+jQ4n4AWFrRQthLxNiJhi5h1JxpN4ytnEx/OQ
pROX2pHca3KoiHDtB15pyF9wTdPPYDiqIuhtSsLn/D0ywpoxRzeCI5DmzdeoKSj2ZlsABaycEehF
woqGiOOm/26LMplW22+7XCwA7HnOwz3fxrucKZ1uv8ficFJ0+joJ0U9g/3VB4AkNJz+C+WuvPbKP
6tCsktzrw8yHFCtqgdZumB+LLk+znqHsf+BIUhtEaLScHKnpESFMaaX5jC5xdwutAbI+Jg4bWwyb
2EQN0eiTPIZRT5fv175OLTHT7AUv5iBGCdiLsRliw71a/fa3CZOpz7oZ/PGXTC6UjIKpyZfWWhRT
Tb1TM2caU6QWLx2sWqbaFJuvHDpGSwB80Kk29b7mspmuvYB+89y1U1qpcsLIzZOXNesJBryBh+nS
lYqGgnsVTHGOs+fpGmaSt9QHq0zYIJCpqf2J/jOZ2KJT0g6y4YTplJiyzhEWDpIBhgJ5eDeJhaE1
Xmh5XDj8wfI1+LWJJ5xQFSR72GYSaN9f87ucFzjB4voYqvWlfmWYDUUyU0RY1L0epgXPBc1hxDut
Bq5igGoAMitlG94tVT5UxWyJRvolkTgBiKUVO+0jwxRfiXXqaqd6kpswwUta0ri8i4Xw5OV3I+Y1
KveB8FwbjBxKS1OGv6zHaiaF6gPm3N2BfDs6X6YlumNV31GFJ1vlc5TcdoY/+s3aVWRdZRNy0bGu
o7dM3/V71yH9Jswq+lu7800Vwe8SKWjVWcfmgx+a8zlOEG8YKqKLuj0ljq1eo6zNTjAh6dgG5FWJ
how1TGp1JIxyiKGxZ7+duXYKIQqwIsCLIYTF9GTD3l4daMigfCzP9cYBN5MLx8YR/wUHBM8wISuI
4dwJjG745A0T9En7lyqIgL0K1WADbbBS/i8fkmmgM8wrjSt9f4MPRuAOnaAdkaX4AW9/vAd/7GsU
pXDAkuqWcWbvMBACUCUSKIhT+ykW95C3T0yu6jk4in9DjirsmvuIlx0hLiLSIcM6AiMPOhLobNdg
efO/txj/Oli2cTDkND699RuBFjLwI/pbPsi7YHg2EOoIe/+M9mrIviCgC0K4imyBYXkVmcR4tMFG
81imlGUid82eoVFMP/6J24kElX65vqH23heAo1L/hWfQ5qtb4QYYswzYy/r4HYOw793HSCg451Wq
DKiRDJhjrDH3m0S8hzCa8Uyj2T5w4JNChPXUoPYNfzdBxjDsnGfxWStwtpITemEDfJE2VHF0mMx6
KtdIQN/VGgqfW8m0pQRsEsAiR9BZ03WsMkGinrdM/du7+u3wN1QPHjRfQJFZc7syPptAeQFVI+Al
nWlsVyblsmRm0fJZPpYWV3EgiB9e+yfNSULNqaFEAbGppRj2K5hAyipRgfwPrS0j+3dS9JBsRLXp
bgqkoucrdBgP1PPmcGMFNTjlJSqe4tQkRjuXLZ6sabCA7qi8PtXC+ZBwaJoGDeVckyybrxLRK44W
LGb6fCCroy4ZFULbooHr1rg8sklcFhNgasyOEjEx89Ybj0kc83TXMjXU8pBgnl2n1zpK4LBlfaVw
fMC01gvahe8haI+FitWsXluLTsFsGgS+NpAoqgRHaIhgvfH8gRcFARRsbH0Hc7TyYGmhIAKAJBnd
4EAYJlX+knkGcFsxAiiQW87Lz2VFGEsMhEP39Ymqim9NTaNGLgWAuTe2oMWk4hKZvqefAzWcdJfr
N+BRDyIv2/e8Yb2f9t3K3R3rPc9RwAveXLwVyabhhIRvriVmNaSa3/e0YKvKeA/mcACtEoBDA4lA
Otf8VlPh1cfoXT7NSNa/vMJ2C0JS0vhjyAzUZrZF7DHaLjXdbbEbeGYdpBFCIjv8MQjtpV4YNBJe
f800+tztASVL9pcUJjopjf/sKFoZv3oB69tMMfWGo4VXNyOwBdkyVsbYU4tKeLQ+Ejq6o8JEKKqt
OEaHuVyQ7k4kJfhwt4qoMQCr+LbAiNejMmkVP+tqIQBvXY4YUAlCKjCd9u6jO+6gWMAqwaiGtQds
8/NJnzg4nR9f4n7ruKG8RtbgaV7ep5ov5RHgSXxa/YHgZFINVyAK+AvxJjLrZu/Yh2+0Qsj6kFEE
9NIiYj20JvcvNhHCqsVZJGFNox+kohQNQa36Ft8mP67fG3sqabg25iZcSTCPkL6oovXsSMgXEN8X
fhtvUgk0zQKZgTjTCzadBAt1lQFZu4XgMXMgwCdrFfxGshKTnHVaUreyY2OBd9MFyGmu3fA8S6my
xfklKgEkrnMrfr80WzNRERo3Dq9sgZ5FzsjsB6epF3jEhLOpa6bzUmKPaJ+BU3ZOLl2p5X+GgaIx
oixIWpprVHuCpmX+/f1ipTzf0yCA+54Bq94IyJ14FJpGlVFIL4An/wv1SdCfR7NLo6/AEeBsSYfs
yx+E3P6rvQaWbFctSxsCwszEYU8SxBGfrxtMpz3j75PWvF359zzUQgak4i0zTTJyP3ZSsC+PBeWs
0u15D7sHPCPEMygN1e8FAAVxFOUkFx4/lZi1spLExc441k9bzDI5SdlQSDT8HqJpfOan0ZEiu1YB
ua/9HHb6pmLcs3BGOFuCMmlrb680VuWjfrQyycjBwAdxllkwbqg3lsaXry6A5yZQMtmXVxB1EdEL
xovO4ImL2WINU0QeJWIjb1q7xfAA+mZl8Yce9ny8tiHgWIzoO/Tn51IDTDPPwxrnC9AV/po3sTxj
NN+M31X4c6Mn2SYn/rEDE7F5BbeWvCK3kncVE42+G4XyU+79dBTQ/7GKafRyXY9oNn/hMhEnAuHv
Qu+v8TDsNnm2RmWA3NTamXgM1prsrg4tSpbXmbWLJxib9MBWWJQSYf59BYMYdz38FwxERSq+4JK2
3ExDKStOXTTEiApw3iQPfWvvHXckBBIB/FeWtRcLI6/Vw1AGVW9P3P+T9YyPd3Yl6fJ+BrXDgd6z
4qU0Ooq6xftGieoKuhh4NaHZeUdIZO2nKwjlSmBmofbYLgeKfKHloiXSAkqtRNASozLbUmTGxNfg
xUHnUOC6lZ1vxbDtj+qVmx0NV3Cpf+d21tfjUY8RHlOsJjGhe12q1ma58mnoUIocDxDqUJ42L5q+
BCNF6pD5xOxpVQYkWj2zO43oYkoiInI7Tswx/cSiuGHO78Z66sq8NxXslfilpXevo+5Cxw+BPk3a
eAh8E+bVj5GmxZGOKpbHIwEfiIpTalhJRfr1lGKWCofZW0pHY2g6NA/A+S9PbcqIXaUn0G8K118P
EPTY+CP6Yp036g1mMC2IzeBTsOqjeJWPatNcB1iFjBlZP+xPtsWk88Mv8ASqz/1FRnr0bSH/Wkan
milw0VXLESiS5x1hqO/F3kdFC5IqRjDedJ3xF1wbJ7RE0sUJOrVsGQvtfRtLAKHujQFKXSRTDx+J
U9fJF3ECGszqwGbCmAPXPGJq5bNX9kh6p/GYUgotDPl26JUZ2GZdQEiGsbKcsS99U47rne3xIe2e
r0JfMzKEcTuoSrLgQPmmNiUtISPAskCr2DNPZcbUXv+iF/p2SgM0bKVPBN9/a9Qy+cZRNQoy5sTl
XjgV3vOCIXNXDwHOddyoE7xZfcxE3lYJ/Rg3EKqPDL9sq8/D0NK8+hgHE2ZAzBMM/53iuokZ6EkO
9ys+MLEVFeoNCiEK1CIw50+/QRWDgo+hktOS5DYu+kAvQNEtWPHKc7N07JpsGZw3LyYXeN5xxXvd
HK4ovxnPUMJxoSjc+NZuT/uDQByxj88+8oNNoL0/wczbNorv1LtkYe/bF1rh/jM/MkjHeGX4l897
abDqmBmKU82yNCGJgKm3XDQSJn6PoYI2n6xAqhV231Z8s6DJVaU27uNxvAfF7U0XRo7xZMgm3Cje
GdYu5voBX+exxyH3NsZfRLBJMjqqRekK3fv42X1r3B8OOJaqqGXKk1sMmW38Yau9+8DT7r0icNYx
AR7teCrJjhZXlrhFSglr8CkCylYrEwuCOp8+lgUHL4KWNLMcfvhAHZ9PQts/c3Vo04jr+mA/oGOb
1wdaJG+iLCsksKLPAdndz9L8IMCTjKiNAw4BQOgJ95BOyqkftAmdSUhSPZhp3q8Jryea969gcJLU
aatITqoFhiaAfep8uaIsrWUkjfOdZSQyEE03taZMDxXRX/LdVj0hQyvYoiyEwjWL1E+x9bt8WVFv
WwK/cVrbyKuy4VXh8WWdACdmjEOjeJqa2+XTJWhNl943Ji6+n5pyk/KthiN6X66Q1vbXmw3bryUo
iKdNjSuFVW2nIUf3CZaoYWp2iTB2cy3fCs/JZ2XX5GEtG5LFjacNXCYQ41oLYsQmewg2shXV49TV
6roDYVYynJQHhZKzxxU/494TpA2s/xwdbG8kIHFKZyT+TlVsQRU8iqbUwnQitueXXf5Kes1UkinZ
A6LWa9cwAo8uAFRo9uEYSrwnli2zTi5mm3WAv3dnR2JOgjA9oTcRgT73Vz1VX2SxLAyLZmXkqud9
uB572k7ngmiMhK/H/FvKlmaTwA8hujod7PvPFYrbAG9SLhcYs5FxilpJKzWHM9BTwrSt6EpdsTG7
OjwR/X1odbR3ExmNVLpk02sBC3MieZRsqx41IiB9RoBX9S6qk2J7kCx8HR35FxJWMhX2hxkYnD5p
u6yF6e+sQWnhktHOssmCYpTqmoKmKYODg4pOGlzFJaEYA4EFCnWv4o1tD8prcu5ohTX89xcyG9n3
rpKbHZ7rv8bLR/OwLoOVQ0w3otDaKWpd+g/DQHdeB3RGAuylw0Caxki9UDPT50zGQ8Jt5tSpCUMp
aRm8b6XorwvBhmMrHmwKSpX4YqT7GThldRlzMlYvWbO2Vyx8s+D/scuTNN1OMpRvOIwFuf6ztqjG
f2981XitgNbqns4kqY3TIO6FyiSM+tQ05o3sotIMR48lN5jWJgitHzH3yp0C8njnrMqnMj12kJul
VAbkaYO8bUDCVbO9fGjiw/sRjCHS0YxuFIUjnBezj5JrPiuSxejbphAX+iCjqMpliaXAjFs4f+Pl
/0T7m/8a6T1tcBj1PHnI6jHSKSAJRKiniKQ43SFxxAdilyjYJ8SWWty4LEhSZNlJUxRDM+raaAPt
BMMWs3yngJcP3rz2tXyJKZnTjX3o3RQldBdn3LzTc0DsjNSeie+BdfibvIAuZAd5GkY7BEmax6t3
dfg3+AihQNxLeFuyryYmORMYuPTUFgF708eoZ1rCWCpB0FJHgiXQPBVQb3m90IoPWLtalvEv1t4u
iIxytz/fL9ftOzZzrBVL3KrLBMpRwMBdr9Cd+Mn2pJDhTt3HPGr3FJNR5WNlOYjZsFrRxUC3pIvd
fPokG5qqiK1Ju5FUje26+3Yx1NMwNehELKuvOR08z7VV+DHXjX8G8SltRjoQ9p96jf3Db2Yj36nI
yUYdtqf87gYkeLmqBv2SzkDIK1PMUOqMP1fuXJSnGqy7gWmRkf39sfxOw7B1nqx5PpFL2YjtTcHf
NOB1M0TJPLjhSFj5VqdlKcUzphjNSJaSYtyIEJYbb6+96Rtumx9/Igq0wXuSecXKq8FZ44z5zuSd
dtY66XyEtsK+zAdz/lWtY0/I6yJ6U17WVqZ5xrEO23On7nTNalOhmI5WIZjpAM+8nRWZBaJmMvv5
FKg5gLuJZxS4+ctHMux5FukZQwg5+/AI4GzsWjjIQT8ALAkEGp7iy6wC7AlTwPCgJewUn4h3FMQl
KcJKdqncbNFzuSpIQubUVgrFoI97CL69O4Evc9DaCK2C83d5nMDkWqKg/Aq+/5Xlr5nTXIm+Tgjd
onvM0n7U057hUTCj6izDv/YocKxnV2DkfJcjZbjuX6NXy8n9epDc+YFQfC8yuMrFe+J3t+qAYir3
6mso6aeNnArr25pohl2lvsKhux61k+Ob83KG/ecLXWFOp9giUHkM3aqS7CrZ/PRF6YIZVl212+Sc
aDP2AnXptVvKwafKduxbIVdTFgYgriE/yk4JBxJtDH3EvI9884iXtfAH/41eeUc4G5xtOftHj5pC
VmgmouERRB92/daloxYfk+adp/ffqr0J7nVDZmpv58fzMv1jGchfImsvtkHvPEWtSMi8LUDzJIiW
5Xouz3l5DH3VYlsAiBhtg+tvtbajO5IPTnucrQAyXiHpo9cpgkjqPH1QRsVWWFnkHxVPzidXaJH5
UD5+pqxG1fHnKndLQpBpnZInAwQfYGtBn7jUrleaMNmQViF2yChxgyOm75UoHUPK2mZerUVYRuRu
oMUcMJk3XsVx796CMFXqNmIglE54Bue8o+Xp56cpD6sWy6YgdXbmGQ0NmIX6mCL0e4pApfx+/Pzh
TFKMHkSBcQivW1nbnBtPibyVgIoxmWRvFqJ3pQNPkNnj9nCASq/ILOIMqy7OV40Ie/Q49Qovps++
q1WM+VuV6atPzNEOzHd+6LC6Do4WcdN0pPwIfXzNHuW7SBGsOMzV8bjGPFQA4OweBCMlArGwPAHW
/OX7f/L3rIkfsepR1MCc3qdJ8KTIXIjj1anqQ1x2QKPBokR6NZZfWJPWQuHTmrTe2ZVdRQxeLh12
a/GQEZfWxc/T1o68gKvr04m6CAHmV8DOqRTDt3nqrYHPTQ9AwlgHRQGBsvZRs6UsX/RKAxpezcul
eFu7kW8hnIYz1Hlw0XlTbLh93vjwskdE/P+XzrgXalIj+bcgSLPf/s7FFhuCGrQ2A9XK4aF7U+q6
FT1WEKQzZULE8MA7gRrQsvUKsJI/bvswEymLSNHoHwEAciecFuVBNc7qDHjV4HwQ7K/Qi/ycvJBD
LUeudOT2H2hAnL1DY8X+H2JZ1CAi1zQMRIvoFck1N7IN1FXC4oeVRML7KB5kN8rageP59dgD5uWt
MQ8Ee+ByS9zj8BdPkEX1L/gCtW+JP3Joo+C48Tu6HkJwTuhpP2XycaR6lJSIQIXIZ28aT4zvZq2o
R7nPci9Ni8SNu2DgiwY4Ucx6AiK57YbUMNQARAHhzF7gQes13ogwhkbrGOMexJ9akmAmKxHbl7qK
5Icdcv3mylofEEOOjGyCJ0Mg8qSXT3qmSPVcsmjP/Qer/02dYMAviC0bJp9vJ4PPK36XRKR6Wphx
ID424LarBQJh6t/9hTbfJ2pcfdR1IPLQQgJ1ftqApN7zK19kL94RCM+JsyYZcCpi0gD+3IyMU3wi
K7sWRPkNZzfnlJ5CtBN+qBY6kogGc9z8RLM+A8Qlhvjk3rHFRcFzEF2i3wt8LcjmIulJvX4QoN8i
yRlSWTU5a2fR4rAyGct7kleoDuk7fTmYvNLNMR/ZaPU0JVyzSnRMwwVN+MwqLQpjYYgHibFbmBP5
XZKsxcZjNsNnwcCpsHUBL5lRZPPLM7jyeP9h/Bw03qSiRkhSj+GpxdTZM5yjhQFuJk1aXWQS0Pug
9/7+V5V+G80qTMSehqlKaCAD8GMfJXzUhXPWhl3QLwplSgiGxws4NkjuT4PNpIrQatuHpX19tKaX
T9ktLbdg+p+HkLVNi2sAq6dQRcVEEE1C4vA1G4v98MuaUuUvkbRqtpIGsPbdQdhrN+FhlmM6y1pC
L1wRwmRHvpLnxo9rqeNUk7BeimowwU/YeWTJst7ReI2jMZOpf31Nrv0TCi8FamZf6PCgpOu88yR/
j/8NV6HZanezJipMQBQuXmCvcByJNUfTf5ZwSKCojs3xOfrJcx1xObHy1PHC4lAHoETkHB6pYk6o
s9VkXg2rOKNzAoHDdAfG+1Q5lxZZ1eKncEulT50ABZYgFdVWIMHEDEbr/Pp4QTGwhM/A6JwBQDL/
q0MU9ZazzstM6uNezL+IhyPUm3mT/oio1pZGRB4JCDzqBjr2ABMFcm/asnTvFm7FlkljJ6gpO/8m
dmj8/GXHqJKdfbS9N166EKnSx1JDuIQNZ0CaDCRYU7sS5UsYFH9YXeq0oux9vUq8ln4aPTcJbEIM
vy7Q/bmQ33+uB10ZKqWqIVtjTVpu8hS1xxpgNIwVredh1QGe8kKfbiCJkt4VgjY67GxS8fnGZ9DA
h38iy7jn0YXh5sxQyRJWbemL2Aq1vfbogPOEGKyHJqClCI2x+M8+RbW6d6wSoR3CFmB8KlW4IULx
s+K1wu84m/KTpi6NeLDyxwjhxxIc9HgdgPJ+p1UcPPXbwHQ4ZO5VeqOSlCt6r8Dix42gaCACYsUR
247uMl1s5AO8LBjphYLnq/WX6rgx+26+NACdmAmZEPN6v7LfSMlFosNlymTRSWSGAB3UdNYplG68
G8qTM5u9cXqQoNqRvb8QcVINRsHkJmqZ/SdsMbi3BfRJBznNngkF+DJYlPo9HXC4WXmXKsHJMPhu
TLQ1WKKkPZVY2fhyLM60bhPiOOvxVe5P64dv8iVKrbo1cIdKb/7hoeT/A+KUO+tErxOUXxtyTp3D
ky6ITh6qi8nXGUO7N1DOAP1JPA4fYJpS2WGM2oxHWZMx2mZsNVk6qJjGVis3JaUlC7MRQdaW1Mkm
L2UUqcyvualaOn8AaKFukNWbA3PPnx7bnmPruEXEtadwDHPEoQYHp7ce9HftfExy/QK3oKx0Dsh8
2PQg3odR3eO/M4j2OYQubhoQGGxBf4khKwRjuf++MdLPP8xv5GxQpyEE773i0pWJiGTrbpRoBzpz
5r1KW0S8WXPE9rcO1jVXGJ/zJ2Q41cezWE6t6yLPBctxussDngirkMdt91sxM4sSRwr5zOZDG+RW
EJHb/iCoMJ32noNdPgIa2/5TW4pHv4hxZospuY26jFSG7brJ4ZOKGtWyXDZmO1uI5dAAyqU3cFat
WCImzEN5EqHFgAvCRIHuIXYmAv9AR7dJmDYTTaAf1HMBsfEd41Z861N7ZAqSurz6yVzpUB5rt6RI
xPAvayCpNpg7+3bV+nLPBi0dB3qssxA6rmmwkZzPQDmAZLFecaEH7DZcgKzuNc7IfpIUhmgc4v1a
YXmoK6Owpma7cyUu/RaoAytVvTV9X5HEgadEwlhOUw6ePx9y3tpqhOAXA1QqVIwmE2YjUdKIKIrs
fl4Yw4d2IqdWex/dcnX5ugVkCGwaF0k2eDV6TACwrDD9uas70YoGDnOXBcLtwnAiSWLbzLIrf6bT
M4n4O5imuCSkJh6zxq/+4Wn1zUPZZRUnyBaNFOYdglFStZ+z4Glil2YcoP5xtalZIDzVprx+71j2
WuWUIMTrhXfljyzH6zsw1/V/p58372EWevSA+weJbZTLgyxFQaILIhW1cIHKlrL5Lf+HQC+TjuSH
wiBfhviZ8xjrrgl1zkzF4rdeZZkHplebKekyYA9vjQ87RcsHxBpRWOXK7PPj3wjzGa1Y5+PaLynx
w+1iFtXJ64S2ROiIInanpqc6n4lazE7R8os/5aRWeqm/uGiWyZ/Zf8ISUIsiuzVQT+fjXdt/7+Ks
rhZtzzl2hrsz6C2T6voAJjIj6kwVIM6mAIYd9SDIwLFgzE3AWHkMupGW6L1wlKbTjE9I36QKepsD
V2Tkre0qv5WrYgluO1nqVw517jLR9uFNzGrCvDv2P/VHKTG70mdTPSQSpRY+kHNqc8NBAEQz5qW6
Ok7jX8ySH7fohXIsKednafe4gzdST+GjzQ58Fq47W6glVo08MC1z0N1B1dpZcgG6E6Vyl/z7v2o7
k9kMP8KTpnfUFm6teSe04M7a/H/dNJSafmHVgk+YIcNso39z7t7pW3vNNwCA5CtMx4cvUby7kS0N
6qPywrht4d3IkdeCuj7FncY3UXyD3GcRcRv73tZ04Xg9bNisfjVz7ZoGxekkMVRu1mmOsYS91Gi1
p12YkCwY56c+T64wlTunZQ8fNvhWrvfxpOl5wp0P/QCNN1IX80hk/SMpuLg30hct4WKSwuBeEhWT
69k3kkp8LTG0B5jSPldR8d2U5qy9Clo3Fug5ki2KqyVPJkVkkc7Xrj612rfqpL1dDe/Dr5LuKlUL
caCKxgsZ0zLGIXrURfTtyrHhBtDTnRkLWlNr0Zs6KPbuX5rlgs6fx8WHM5mt4SQevFkkDAiws1NZ
5PtztLqFsT5Dzt8Tryio7rFhCOsBtn7m4Uqi/t0DsxFb5ixTEk7De6PUDEfWlcyO48QsngLUHUbR
KvWMGX5/aGkG4Bo2wsfeJKHCmFQyk0jhZiHYR+qYCZWubFb6+KKpUgLCPA6l1KhpqaBIKBmNztEk
PnjI4+u8GOsRSFfMSnDPZVIrU67dSZHqN0cXaRiihjJRmvwPd7y2DldjxeG9r9C5hYxSUgkMnzxq
nbSdK0NZ5bzRoIbA88TEZ7PuRn00asvPf77gMsamIont6GMOQSt0ZKmxbAweY0cBVSgkJacjb6KD
aCpkbqFeSPl66obaFtd4gwUVQnke5fhs93ehgSkiqmvZ6WAUAR5dc3623JYh7/355shBO1xsYb82
rcQcQscv9TZKW7wYKQ8wenNU26IdRC1rtolE6j2ZfYBuJJAiKb6VZB+Fql+4g6go0ZPlEWCKlURg
4yULGQ+dR75cTEEqtIOAuQSeS1J8wDCMYOHjGHQkP+Ai9zCEto5d27DhhotCWUQ2NJMIboLzyLzb
tgl/+lnttuxSCDspzFHrhLSVQHqtVAsMnJcrOIQQOMxCvimubb0JPbCPEzUKT10BbKx+d3ktAKHV
CnrxkW60PFXRtyvtCYlJf5OrUAMUpYfVRP5bvPfjZWgg7c79d2LCebOIKNQ40wb1b8ercZGwRcVl
PT1mTFpKdCkN9UmvqFPyPPSBf8+T1QwrIWFVKBiYNZskbDAxnl6pHQ8Nz2CjKiWbAR71JaR09bHX
LggY06HQkzkEpYiCaHvbipnwhoWNBr8Gt+EgRxkowX1xa9gmw6V0Ntlf5FGbFhne+3kSG1h0NExO
98UFL/EgZKLL4ObqjqgZVEUGf8S2b0sl90mnRZOnI/qvODaLxxFFxVZvGDkF5gXuMT7PyMyhh9qi
BUlMr6I1yuyRWfxK1LQGJ196OoNMj3icfKs6ZLo++akba52QaLp5HK7IEiv5Dgp32UJT6DlLUHNJ
orPYZTV55D068VPHzFsfAf4x4ui+TS7PucWJbzHHiwFz7EfEbTdBXS5Cc4yLYFqYpd3MXROkL7Ng
ZJldZx+l7Z1IpwG2yBMSySpdIgMG4hdOJarfNbL33t1+3NXpZdzCYvrvl7heD3ygiycM5i7KFhJL
3fiOn2RZDTNmB5gby53rghscRVKnsLnU+Ti/IUvaWJ9uauwXaMSIwYp+Rc3dw5tv26Wz70J0bWuq
yhl6p+IbufPc1VoxNcvNpQaePPs56cANcwSSMRwxG+NF7LjubWXVMpvD5IIs/6mhSLCZQ70oq6y8
0VkXvU4enH03LftkXf2yFrwDpBPhYfk4SxfCi7/fhHXehnkEuGP2ZB8DZ5NegcirttN2u4bFrRFQ
lFfed66WvOH1aIzQdbzJX24qiDixn2IU/k2hMNfq0JhZ+wDE+9WPmBz1PwhQzWDnjyFBw2l/q9eR
9WyHRb4119V/fwikmLHr768uBDn59kOHn4kFbZ6k/WoMpghBB/73g2bKKVVgEytMUBRuiHBfNkbk
v6D/15zI7SF/Fvn6mTC2C/mQgmxqIgbytCBKHjKDbKYK+PU5bTbNyJovKebUl5KPaiAVvz+ThwEs
jIuVllGg/kETH3EL/OO2tEs3KruUsNL00wp628BQx5iVWuFXFUzy0wc9JbjTFudc4HKVdXKXQshR
/sKGUmOLhhZl7oOHzf10aymJtuokMd5VPt5ZA6VWK+ppFrBQ4Vm01sFOlupTpYr+EY7b9q6CjSJQ
TACNpsvSXVBgVs+gNrIOVXRTpU8PcMzIZRfiSnsLLV83SX8KA/EBMkJAL+B6V3Len9O1x00lFDmc
+0fo7TYMoINtx6uN5YDN4tKFHnAuUPRrG4yDmiySMAfWqlFvQSzYfDKdndVBlPBejz+/kBKobsQc
797rt/oXRLLrCLktN3d/1ObwITB1BDzIZyjT0Euah442EulXgJNOkZjhSBGykVWCaU7D5CG40jr+
yjFMFVxzi8t2+jPjkkdifkjllOQ8PnbQ31OT+7hdBnEjfYGYGuCXCd6AH59/9NLQyZe3HbJIM/XZ
ePJUmZ/caw6DRMJ4o15TehWLdw9BE28uK6+DXD6KCSc2pDj1HuvDqjGmE0OuC7ecRD4DEyzQgIKn
/Z7b7+5iBewa7fG01GgRdE2kkV7sHPMzectPNlcdrsU7xmM07neDEReIySr6w5pM/XD2qCmN112/
n/XXYx2KpUlpA3AiAXeVLVjasKdUpJ/TGA5P3ihdlBNInwyhO5O7xh0W4eDFx+ZLbLHjSW8VxSJr
YMtN+/oKDSqfF1wcCEovNSUh/YoH948UBw6V5pZtQ0XR9ltUQ3VYApy5mupc1kdwwPYSrvkAOS/I
WOk+KvkMQq5de0hD5wFNBAIdUYnWdrB8yGY0LSVtPFv6eIz6wHa60ILzCidD+pS9AKIkAc5c1EkR
7dVXQVOheR8k4k/7a92+4qaBzZw00ffMplNdpLgyuRsuFVlq67Il98kxF/WilgMMesB+1+zb4uVu
BKQcg2TTmiRbTMYTgyDRn10yDrDj9RX1719r526lcKnQSFXp5YBwIVviPXPyV/txmzwI7/1TOOtH
XXIUCO4qZiTB/9m1Oe+LFemDHSA252BW+jQVBHomqMRfsQ5vUJVK3SsNfCy0vOU4C7mWQYNLApE3
mlWYtHKMzJRRsNhZy3jQzOERPQUmQrNVYlokXEpAaiF/QhBXEJ5jqSh/8k2RCd+m/y9IYGvtLx8Y
Ko7BOZcsVqmLqOutpIvBCF7+MLOP6LSfTCO/hwQCz7sUSUJSHfBjZttYQBNT8n23+DRHJNOPQdph
KpCbzpoFiWoal5uzG1IfI8Fod3EiLdEMZnI12eom0ZEuSrugpHPFLYJQKfUawn4M8i3rfgaNY7Io
xOSbMxCuzHwh4UlINct6b7mjUglxaPas6PQsWvnP3X2NMVk8kvuJghUiVehHYQd6QQMD30U+lO4x
3xahoTBmHGShZDsuo36iuGoN/sTtKaHW2rLDFvy4+/x+bZAtj69SUfd+ojoNj5AzSquYcDi5+ssD
Xpoqi6v0TUhy66I8W8U5TOV++rBpn+gc6JSP+K2QlK7SeLv/Dg2buiD9E+fQinMc8FPKgWiSyt4v
lvnBl/ZD4DH14PM+XM/OANE69AJtf/3F9gKmM563H0c111OobiGJtuQu9whjrvnF2OLti80WSqxZ
ll6rHUlP5/DTVpe47ixe79SXFPlAzE19uoTBEOHXjLvx2zTsrvFUcwfPdtE2uOjgmU6FNlT+6KEB
7+ZTPQ/TO4vEfEu5/f0OzLwP/SOOXDhltSAjZAmOTDBpgkWld2UcPthLzBFj9wbZgLQ8lV6eP3By
3Li/iBu8ZXZ6APjqJeZ2yDkOzskZi2WLe778XH/KXiAlhRA6nES8dskVThkHcyOT2ESgz9okgg7t
mHwBlk4UmyCdJG+jKvjxjcIQpD3f+tzVENtBDWO5CHNjoH97aJrkPKdOU9RaePkJKOTpBn2wdUmn
2jzxGOVQ8z2gD0e/9ktUkFxIZvy08qTinpOIoGXPS9RoWkn5Y8MKIX/cVE0d8xy3ZUy4BK+94D33
QhldjGRHn2rejBCN02fntSzSSRIPA1U5n55l3HfjHi8s+C5cpetQlxdPD/lxJNaznNDyVXa1/QXe
6HOlKq8/J/xJXM2uG4xdo+Hz3gEHCbxvYeAk70qNLc3PcZwuptRlKLz6EiVY6RbWcPA7Goz7Gwgx
0YtNzdL32ez3BysVhDJ8Z3vphoiqXFp3u/Er4+86uBZjDTAdecEqg2ItYVTXCH01uPtAS8BvJalg
M/Vuu9JkR6XZKCNNIJU2U7OUMYAGs+HuimkpZd61bZNSRyTHPsU1/u4Yp1EZezFffKHBl+1yBxv6
G+Pydh8hklOq/+Hzv37weD3eByz5W2pZye6RVOADBI5ddxmXBfFL/oAa5KYy+FBBIljf95qbm8eS
sb78VEiWkqJX3tr1dWcnmDtjTT3sXpwmkoHteltwy8glBp91oG0AkZfLL3D/B4JJ2SKx0oqCk4wI
YnrwGZnn1/kTN/i/tgIWYymt2n+fVVtCrlHETRGYIr3MlAd60xpblFYfU1gcJRnSuOHB6+BTX86m
0BYDV7k1UNf/2S9/zBydT2hIvuZ+9X4oBhPbTr7h7JglvWQl6JzTKP6Ufb57y4GjmtM3nvrtKQui
wcq58gsRTdDwvoPwyA801FnvB3S/9s4DzTw+v+hMLgtc63On4V6E98ypUS4yt/gktnluYtMUbqYi
LSZSa96FROgh+t9tr6x3PAjM5DY83CbFdDP7WdbjEcVpd9X0tXWOhSNtIArotk8haGzrwKa8IuHQ
mZNs//VGwWrTntckwknmm7rdj02NfaR6aVYgm/hCA857qhYfUYBHgGgCJsL55w+uZEMc6iuM+pfo
SsLmU2jizkSEDs/I3jLKkWPneqScjTI6+GmvxaX4E/BCCv+tq91HYV63R7UsJUytgMn/mxhcYpk2
B4JGed8damssEGhIpZaJKia7BBUc79xaQC60H68LzC1X4Vz2Mto+GmvT2jVUVe9geexBzQ1vNfAK
IlXCmnTL77C6hf2JC2pNpkPfFd2zmO6Kb9hajiqeocpAkqFtE5Sm+IhpntnCWzf6DiNNdbOKhY1F
KtJjPUPHEB4EHTZUgEcnA9rHdoIEegkcK0rnNUOqFZFkWUL+OgkGf7rxlDQYYZWWWRD6byFtaQ7R
ZW0rVocyMbIdl4/prJsM4ACUwrfIU54K3XxT+nvHFEKIAx6J3GqACEctkH4w6NCy4HHmYvMgM4Xf
0iFO8nby6PmBjsj1unntbO68NZ6dTtHRGtSGF82lph4ydBpGbRke9ciZiEpSYwBQfFUmCWI2xhxV
PZD1e4Gyiv3FKbT1gkQ7J6BPUYu66stTxKrEeZ2xnb0RfG0Z6ddteGnub6y11dl2ETh6Py+tF9Y0
b5Opx50FU8GvGrT56o+xfagxnvEj9Y11RvocXqy9i0GzysYhCQD6cddNBAp/m8Z7OR3INz0pSF6R
wSX+ASkKm2QrFN5k9btpIBohW/i3u+ftnT/n+NVZ0cMd6jEi1sJGrwH7nHjNRrmq6vSPpT+5JIre
7UQX4vZLBIVWk4up2vh2XrRdYGcXa2qrXN7f9YpnQ6/63xD/aKBskhGFgkPP9O1bGr6E0MNFsgko
Q0W9T27byyjUnbJuVsBMpHIA/42iqE8tY4FBOe2izrmHYfDMIMYc1e3cqvFtkvIC4XFoxKw74vA2
z4q4kq0RhfuZfwdEENNXkWVQojZUctLc1I2j7pTnSyp4JW4U2u1pvpRjwAYyA4hwhz3pqbYuFm4h
T5XPD8G1qq30AkwTm3+ot9luIPE3Oh2hc/J9JCivlslbVk1Ff2GK3aDw+oTtCuiHt/FHeH+uKhRg
KIt1M/vLaJ2ZuOjpmOW/wptGSN/9Xp6uWbdqWyz0SbegetpOsOtNuKWCg05rC4998q//cIacu0d5
ihMxAne4tzYAfIbvVARuAua24nlGk7mvze1X2Vkcmq8AycKvV/a4m6oEQiRjCvAovubGMxx0ETOP
6vkIemZzgBXJLQIfT7F3e13RoHbUbh/EKeCpM4Aqt22lyDl4jcMLRKpYxcn5quyOmsj5Zli51ldD
a6zYrhGiGrWPChzYovteo2Dz/BEdgjdpmRlcDcFVPQGmh74+l/bSvQvwJc0CVtn9jAzNX+TQWLuL
5G+/cr/71bgMbYi8Xq21+vYiPYRVo3ITbuLilwhvbAQpp0nGhufLwcqA0b2X9mwDFVBGGtwJEtfR
dSKmGK0ceKtP58RplFzpW3MIQxSDRy+9xy1w7c0z7seTbE9R6TZlRLe10K0ABOZ8pVCET4NC8Hk+
SOTFts1RF6QBlsyfjQAgeW3Y0Q8NIRq8JGQf2KTWrAJuzjcyUM2F7CC812oGyIvYASbWbW2Mvgaj
68q5KT6QzXmLmQoWyf3CivKPIzVupqlLrRI+arrnnNOdKkV8geKlwri0swt2/++voVWf47sirKuL
ITnKDImtPV9SdvY7lKu97dCQphYpHAtw3Ft6NbcxBGpA6b7LzATkawq4z+glaW3Aa9oDBXtWNXDB
jljBXhleBIXdWi7QNgfhRmPJVPq+5sy6BfAYWP0HSkR9AMx9qqldHAmWeZe1p8EyM2TDaG0z4uCP
jafAeK3BbBfwmtSRTYGMJJhJ3TtwqYxJU+W9U60mfV/C9yUes4EI52FP4OcVBHTp/USBqbLj1m6j
TUbLyhsfcJBaP8OV54tqatWgKkePGmjeJiiolqbjA+PFr5xt4WJrp5tx0lnPzUQ312YFMq3wUvkT
gDfp488Bi7dR8Q4a+DWbmsItPY1n9Mz6xJCbEcRlEOqH++sbgSkV5lJDrFjJmmK/FfiYqHezM2fy
b82rN4Gg+4qhZeCuggEe9KLBklmJPfNox1TAWzmmvT6J2SO/3EfviMKTgS5DbdWoWxnNzuJXTu6P
ACsT/Gt0oV2s0zeVBalTgpyyYVclQSrY+BIQUL45Pu6AfhFtJg7Hj/9k+AvYoTsEI3Bw8wZdtSnO
ReSopE2GjkQv6Y4nN50dGLiUB4hXUZVLOME+17iL0jv4F0QVugyGitpmkb0tmlXXRvranJ8NMxI3
YgxQ00paQ3eOQ6CSaa+8Jm1vgh3/QtgdTWnIrk4exWkIKMejZjG9gRrLAjoErf/EHuJg7xlrGabY
ROgn8vCt09kNCEoKAK2wK908QoTwInN55gcukTBAnrWF+UT0frrfmA74mugwxEFYx4oKmJBdQ+OF
YCP2n3cHG5ryc+DBrLnzVYN8wx3l3t29gcfXIR3STwdrBpakgxo7NUBXW0QYBkzSVDiDacCgoyMh
HRIySZ2j74XElKXBj0Th0YR6xAdf8QLG5iNsAqS3W5AzNUY7m+PmJJXc12/oz+v/6kSi3/iAClTp
h3SMoqvZ4Kf+pVtFwCx1Bvt7eE3IlEFFZdyjl5+orhsTs6E6CKQrJhzZsuczKgnfkDhUJKb114k9
oWnO2yJBn3m/OI32rlmMbVDmTaZCmMYRNk9RTNzzTzK1Slq+0uhqAxpYRCzG1kcoZACkVz2qIJ8Z
Cvd8EPAgJPtWTHKQYp7o8PKWYadHMlGafBm79NCcbnu5XOeD+6bHJeY6G7N1pKFi/BippgfyaFZe
eaidX7HnSe3p0komjyxF0vTrjo2sSj9xdI5UOZ6OizRmMfCWUiZ2Q9PdjL1r289HWLjGVNWzZ6Yn
ai3kDeoCib5LexNWeem4pXh+89QOzUAny3YVrZd1iCukOZ47uUqyi0i5q6zAywup2npded5V9NVH
wkrjihiL1GJ4qIGA7wFvCsQ3oaqETsXGOoqQb99AOBtMFBYIIzXgA4SXaM0N6sdns3X0rhDIbRWW
p77xlr8GfQfuduSzeOwb43aaEBPnpzQEUj9eL4yXVvBULnMKhD8FveIZENaqm1UHsC28Qnn98u8m
nyA3A4oXiV0wakwPelJNuVq5RoCIpFfI5KGVGQgYg8sC+pAQYhQybAIDg+JFTsPVHT77mNt+Zf06
1AA5UF/H4yfkkdqqi6VvbzVqbnoJlME6eoheFG3op4HUpQNaGS03eFtRN0uW0ydDFARZtWdhQgip
DF+lgpr/isiS+1tMLh5dEit+OCt4U9GNG4IESb87PtkmK2qF2j06VPv27CleSOGMN5W8kUgvW12T
bQTBuzbrsWRIoOutAmFNEVquqhYZlGNc1MipWZ/kWyfBJSZ2Rf4l51iDsvGm3FgJQrGcBBDpZhqS
563nOLFTHJraBgTd/VJvnenK6dumRwZjxI6J9BUmJwK7ldokd56M2W3rsTR1LQ/BpMrfJHqWKswL
BIv0KrwW1+PgRMT/pbumTe1v0DW2x6DhMRbTd1yuKWqLorKDUCoZgxE69PUkSgCPBSrQDA+KPDDu
iNqqDBP4lBsocQUqJL8r03PVsdn8/nXkMlpmX3rv5pyqlMZgaDNjtFE5TV4HzlhMZY37Q+FUfjmj
PSAK/9+r7ScxsGipkCjW1t9nGJoPn2H5OdVRDHjptDVn0tRWYgOZfirUP+RGMjks3iIhf8f/ZThb
u8olVGTxzF5yFit1b1fe1S6TUtB2SK8OPeBzZnC0FkP5r1/CeIseZsyDdDbYInQVeKpyRmzCffVZ
htq8FrZgtk/cx7ogyX8XeyTwRw1GBWvUc4YgYTGMFNwzxFkyXu+TGLQi787PJomaXsP/AqKbaIDK
IeAb6M1zsdUOCjHUz9KA73c9GawAEQq2amdMbeAuhLrQH06dONWT3ujaOMNwyaADM+8ZCEPtIhE8
ensALitY43sE//8/Y8Kp7Uh1iImYysCfn+Aa+AqO844RlM+Sa8jQGrNtV/3OuE3/2qLkIWWjLccm
WkQhek6vu8GKpPCSNF1INk5Ah+ob9Lv2rfp1S6PZl2CFfTyL3HE+2U9d71QyMCGotCisztsce8MW
YzLNMg+eZNhPx80GYKqE0qEA34F5WLarwEUvgMMU/XP/R88wd6LAw7l20nOsLu+/zlwMjoxjo7v3
CJa0IZzV6lvALFA3v//KiEpdL2tTB9zgUsJhL84L/KgVsWxB22sQCXZdZMsYWe235JPcT0ua6//c
Rxbt+cW2oGiyUTVaibmBxZA9G8zfk3ndnkXtP7O+2TdEbBZGHjkUco5itxUGgp1ooYD2GsV7ptZn
iFnzDvMLw+bZqdXRJJLTVsG9M1Gqj8X2xawTn7uw4PsXymw2d3a1bTpxcaB8M2bjbLjtv/YweC1X
6SfXcqNaS/YjJjVs5pdLo/1YAW9kECAQvyZUwh9vc3DMLztQIPdzLSaIt1NT9EPW0ye+ZNhIHIyt
kiYOpw2aMEI5gnQt1fX8AWpEV1IhXrqswOHl2LaW6GJcm+zMRtH4G/cOhOb6aQZr9ecLxfjI/RHh
7DQ6Ny57/ROshjRCuaP0XZ4Gj1Bn4Zgc16DzUfNUJCWUb3EXOBgR/DW3mMFXxKGK8SWOMcr+e7+U
qsNfIo9sWlBxaALVqtS1QUw7kL/JlTuZ9NhtY8gh1n1Fm1gYag5lEw56MICB5RpK39hNaAq+tJtZ
L69qunzom5Ta+qkYBkUF/ccGsvs70Vt/r6B4fi/XVlg4cqoZtYsvhwXwLBFVP7JeNSsELRvPS0On
STyO+8sj3BjF0/6x29DPQv6P+Sfv7IjswsCQNXwnPpszUAyR9l++ctzQvhrpi84JXox+fKPHdW6Q
byPjLB2sqoj/ffpUzwnccnlUoAswsZcSbMt18ci/vUA9rj1Pvrt1VrLPMZ+Irj86ozR7k9KEKl4u
3jeoFJiSmuuYgPqjkrOtvkmGKZk9xh/z/MORTcavy51lC9yc+gd8fw9RXEbadCy4cGQYx5OvYybD
LT5bZlT2xOvhjHbyZecXvqiWBBxKV2Cfz7vdyty9P8wa/67Ib8wPf2XaEOUngW+KQGB2QJ32z1fX
kMYJeSpR1BCEkXRF2LEP/64ngvbTsURQ6ZvzCnhw49PjXsVLxCSksh2J2nlE9K5JXBhpCMX8rEG9
aESzT2oYgsG5Mo4xr4crfGn+kduWTp/zIWcdF5osHezowIltcs/vWVGScL3kZcYByBQXmDi2zeRz
eoNTNmsyt9/v3zl1xMQyxWEP3STAdDjVeDnHWPb4d+Tfj7I9cppPmqHnhdxSBV0ExN+81Tuq/WG9
vIKgT7d/d4rhPJkD6266XK32a4o6Mbpo6jtgNQu8gnl/iWONXXJ2oDsr75zSoQLN4N2nOUJLHJo0
aTAInFk5IjKEadFaVjNKKcRIHNlm9qx3C1fKNmTD2wCWuw/X/2MCw+sHOCuCNJQbr3jOXb1xUrey
IAcCw+vcOtGRNQY/zsW7sQf1Od8Ez/qrhd0hlCTI1Dd1XiFJfUKj1fssaLdw11XE96Oc0KTrbV7L
Xx9r/GMySZ/kw5txgKa4chF9IqXxAdu4WRtNbDdxNIYXgP04jWMrgrHvT/zlUDUD5HcAxejnz7nB
UN3LqgehMjDMPfcO6bTJ90Zqx7/6rjmM7kRvrZgOAe79A0zx18WaQFMSG90WxCEL552AguOgNyVM
0NMMneGg4xbAhli+oqnKicvw+qBAIoONlqnTv17i4WOHUKmjlbZC50Y1Utw+1pky0rGxz8UNQ9+i
Jog7cMTXmowbv/zq3uKcnuqCWM+xv3RY/AeMW1mf12rgLE9oSihfA9RenqXbN/GyD+vx8UUgnCp6
Ya2N/ZdmfLVeZo+04eY86TqntTV3kUlpg+14qwtAfYojwenYR0pFxTLN90cO2Ju5yPFueuFCOjAD
6YXWdgmFBZD+7pjX+sMJpaeF6NvKYSO772TC3Kpo0hUrOByQr30Xa80wgq4pSMto7jiPjvr4rY9o
hI1YI0DyEERAhfQAtij6zIeVWZ9yvnV20hQz2se9fERrp0pf/VA2oARP+4yCmpK1U+OaAw59Ub1T
SNsmj0gcpVONVs/fNGSu6L6Gke4z6GRuxi9wm4UBoMyBACwSeTAK+aSpwY5/A/j093Y/8hXAtZo/
qyX0AOiYsb2wlmF0t1u/OQzRhS0d0sFK7WxrxM5F9P5TrkSnKRCnqB5LMQJFj050JZt8cKPLFdWJ
WL70o4DY2suEq8sWpUOCQC+rjdtjwj0aPin+yG73Tk6EaapzwbXgV/xrpiAT5pVm5W3gAPFAVM59
DMFBrrG88t4SusMZIZL4l7EIrl1zmhNHfb5eyeGfYM10ZsbGvIAObz59q++q66TiJDIXIc5qMR4W
ZeE8b2RIFkp+w9qDXybiGrLvWeCz5Ow6w8IS0ObRhyp/A7kvv4ksqYQu9jNe4Kn0lFalOFDXjL0n
K4lYMh34T4mOzE6kZ4/ZqWVFZ6i7PlBCFHXHP+G/CZ2CjoGyPi8PGNI0ZZ4i984Bn8LV9gOI971N
FXs0jerNHk5prs6joR0qT36B4S0WOI3/ksVr1zcOZCN5VjQVc/idZT2pKCBH8B/RLlD4v7UcZfrX
3Zn/ibnb86mL5f71cldc/WhAePzn58XrQYaawSCOBC6lIBgMfdyHUZVR5rGHWg24x4pc+uOb1JZQ
Pm2qodjFsI7C7xURNnv53dTlNp6KFVd9vdduo9yC0mjlXo1jxc/V/YnDLo2uCMv+iuHUqanzhWS+
zNT3LBk7HVZ8X9IJVXXLyRP5sgn5QA3n7p5xIoGcDJw8vedJvNbB+H6ke42B3bfeHSJQl1sj8XTv
3xwXwSDU8bGFmseeRezSW9VwEpXIXQbqda52nPZjMQL0gpVaaZ4goQ7dBpOf1kZ64r2K71uKKpxR
NrGN6Fzt137WfpobtV2F4gTLTQr2m6IxyKEAVP/G4xxd3iAUqqvDcZBSjhyvQmJN41ioK2S1xqEl
rjAVyyd71kx3wbrJHzDhvaX5u2FSxBPIeemad+C1XTDv/kxPaYVM2hAR4Px/bD/rDQx1kiamFWvn
nxnbAbx1ZESGIYIo3HDf3SPfGb2HCSrKu0QrfsIqZMbhcEorUr8Iz9Obm4gCmS/UzjuE2C+axxLb
Bybri75rw/Hb4u4vF7WXH5eOfmGLk1Otj1Mymbm8BmJQO53JEUczxI5TvxMeM7laPVDPnBYzenuh
nnomTQJSRSP7ScK8HmKYu5WhTNwwyC4fzU1Lt5ZVn11fhqHx4lfWaTF5X6mo+x6r57Hy101/LZdh
K6mo0QuQDordnjzwUDA3TguI7JkI1lPwmzb1OOR+PppWVWKgBRZB27ucGFEXA9twa4tRWL7/GW8x
plWq+9Q7t2JLQgMRR1l2vzzqxCY+XjRAbdzY/ieoUMjC+M2UthOVQIVSh70mWDKQP818mvYUbvJ9
1efBDBGoULgapITQaCJtr9dpQBTWAvl1hJ5u4ZPfCfqZYSNcn/gvwiy8yze9sP1hCK9AnrH+C0Z3
whu4LCj+4IGgyYF0oJzYNsbMlIDFOB8Y7jp+xH++tQ9U1hCqqogBH4Xh04HljfAK2ozi7Q3WMqhU
9c3iEun0Y4L2PM0lji7yh68HRRis4q2wa91+DsNc1ycyCl0GIZVzFUBcJcbMGzI5VQHeKobmuoWx
r0fpV01a6V+L3hqLgNXD7rZwhGQsEcA8AqK9PFesHRBa8KCocvugjfNgpbvr1ZzX+nzdP7X27pW5
EZo+UNjr1WcdYGUVmRLmZDfeMmNaOh98bm4AbUVKOTnQAUn062BefAp6DuPyOcAx8QI9/9dCw0Fy
6clyDU7xMAFuVzjvW4u7Gb+xwekxPBBo/KH8/ilcWSmEtaOGFf6i0eWoVdNvQAJGVoxtyqvIzuB7
1+4Ou0AFda4iPJaGreei4/3mEhZ+GhiBfcnBKw4KXWwKaCf+KkW+up1nLlIZmehl2XXPjQmotGKi
DGxqX0AZkPPUK3jpBXMRW6nvu+5n4I39EUGYMPepEFvVwzmAwm8lcj5vCVW/Inpp74YnpknpiEsL
HuCa+90b9DyV/DVnHIxrxhE4Mk+NeiuwlJ8E6HNINgaoeKzBeBjSo6+5TOCcbRFXd/Ah/SvFOhqM
FWNsMrLiQsDxjnPX2ENYKzTlIWj4dqAET/uTrFwSDwzU0XVt4cQ5KbfTfwT9jvqtVCja4o9SOwfs
RomO18sIfWN40IbPmxeOMojvsc9GQRr/U3xIHkdVdGJXdg4YTF33vvevUAvRbCpQupDIUoiOzQ1m
P0AAPLKsgmEVmkZNwW3MDi6qTVfa2hYNNS5XzBrMxQPU1P/RT7JdB/CF5/GziCK1Wx3Xh+31XV8t
rOMma7CHIf6TxHi2tCa4qnhihIpzvrUI6F9NrKrUJeHRhfxsmUmFRstwofdRVMaNNLuYFxa64dLj
cgAU1zizsyHGoWr6RqZYe5HkXesJHBhpO6HO75qnqJlFbG1VKYKzgt06gWUOY8wzq3xzyrTjFBaG
FN3mfavnQ/kXBX6erkoWVP5xwXpJsXNY58o4kH0wm8NQg/mopu+1G2Vt1IjyKS9BJ2PoefY1KyPH
xKruwDj/VNFzFjCj+xhQLIbEF6ircTV0gkgbBW76TTATlVICHVatiH/cKuV9QCEm7g3gz+ByisrI
PVmYwX6QxqkG5JSLXsLnR8GKDLJv9FbIlwWYWEqgwpVUumquReo7ZNL1pFYxOzNUgtzaxwuoGXnu
UG1HSSJClmHOQRKbqtYZQTtOepz2p/mAiabmIx6lJPF85T5IDJCbN7lGgOv5Z9abOdXhAwDw4k9O
uZQrgl8s3uEdz7MNbG25gOejaxQEmp7mJiM5VpsWwsuozwYPvMU47mZh+4JvQTy5T6nakH9jMHqn
GmYTCSH5DNq6FaA1hUgJqBsMT80ZlQyNpqHdwGawzM05CCnvTI/7LWMTQr21qzMaezvHGKUEniWq
TvauS97Mx7BtYLkaslNImJX644lk4K9d4BOEBNCq52ZVSneqZIJsQoGXpys6pG1hn3GuWobR6eCD
rBMiOSrpLjTfi+tqV75OG/SoOWF2xclUgEKkBnP0/kWAQXJyQzWfkmzPtmWvEckgQsm767651Zxf
UhMBJL5lLOZutybgKvYWzN7HBO1OFppCn1If9NUhK9CHKqI1ZZJTmePp4yr8Y8uo0LWkvtQuBL25
kQrcR54lhO1a82at5bFz+gWPrdr9FES+awW05d3NMuhYvJehfBEPNk1eemssaRd0D9HOK7xwr29x
/K9JFVbyafTnFZmP2uWZnFv7gkseFLLufSjuvWFXjpHiyxqzD0HPqesgUTvXEAEqP28H7PuL0TRs
O4GvvdcD0mu1PbvyaUD6D05aZ5wcDF6gjU7+OU2+7WbvFewSsMmf+w7f8heXmLfYvhd76zniQcPo
DCoyejPB4EmIWOP0WwrksbJvhqOu25bbRdmetA9L5kYr6FYlrQWUHOx2/eVbXe1BFjG2FbxLkZPa
ka4det+TJ0kTkRrJVxJ4PCsEiakfSBx1scRFyhUwUH4RHHRm4S0ISdlcTn3yrSeOlNinB7wuW1Y1
p3mm1nuEggjt0d10LCl8UMzWOXrbV8dFiFOel5Z8pynQYE2aJj+VGzye/oJ2XxkHN0Sc12ff3kkT
Ra4J4eJR22y2WdlmJgFPgeknDyXmNp0lxWfGq6hwWedOdDTSyczDyc252BIyTDWd+TNgubTOcY/P
rDK6/ZFcEJyYkyVLb/NNCRpaERimoknX7lU+LkC15lcr+rEl5thmlo9jJwRMZif7oW9e/u0kMnIn
HMw173SFNHIcgPWmbn3vfy/mZ/plxkQT07lEYFAIrtf3j7dQODnw+Buka2PIs0WnmKMb3xr0jwHh
YLYzLBgyNJv76VUpDxc9LPPBH1HYjo6V3DOKKqYwXtKGu3OD0p6JE1qsYg2kOg/petlIFB6sakJK
2p6+x++xuMNNOwceuJc5UYBLv/rcklr/8qrIhiDwDch1R9Q+L2gdPt8w7InhTE5HUp4yoCOxFpsw
B7aEjfOJmRlFt4I/R4pE9IoevCxHIorx3memL2p9DcT/VNHPYlRvk99PmGM/6eTozr6hzcfcOeRn
Gv454CSVLDbcpD3rn6Vp5zgZn837CRXhpRoSdTyBKThCDnJU4mwatV/P/TU2jwdzJ5hYryMhk4Wm
XzKXNgui4l/2z6bujSQP5NdxGsuWaxx9+sfxYGNU6CbDu9aBHWlxjnAFW0oeZHzNItBpkUP8jBp4
n3bq8oDiIDhgubod1vehuM6NQB5vHLTfoAEcsAaAy00ovEk7+hp2hN4kYsS5pTqGT6Kbqxsn7sS6
CgflVWUAP6mNKZ2NMtNyCYaRna120RCx7VPheMr5luYGg6tm397BLv6dc8ZgYeVo01kLR8zdMoMZ
5ae8KSkKdZq2TrP2a2U7GloHt5I3PwYPFBqeC0W01vxCAYVMMr4it/0BLeSR6MLk+xqyV75X/ZjQ
nCYe7TAwM0FJPo3IX4AT76a6XPGyRj2egp/NnbF3cKBoUzsyVXzAYn50YQvPyFku8AyMjXmFoNu1
lvGecYl7cJtS0UoZ4kjM33VCsbcRC2aGDKJTugflerNzuzlJ2HFYdHkdkPpSKmu7qs/aSWpXmrfV
mkdI0Dtt/8krkCfbh7gUSjD4rzRxl26iW4zbRorOPV2m067bTprZluLmn0ulqmQpfUIcYlH8TEqs
qlscpx1kXHF/IyUcD2qGwqCZMjfDOmDG18UKVFInB6ArAxPvIsP6Q1AG9juj6ZMruPtVW20GrC4S
tMnWIq0xlvoO23iYE/nQKely4s8VAgsFo3LbqNE6fENOz0NjJMlpvIRc0j7VlSk12fudyZXOoWa1
zOtNpJbMpwP4I3D6dnFLxVoQ4wBgWNXktbxBseuMczy46Li32AIvbIoaW+yiQWK7xIONWjKN1/Ji
CqnYkRoMMzv1oHK3xyOWKra9Tlxp73XUkLSMOGdMvm5WJg9KhXjexW4Lwz0GHnWqxr4xiyBNJ7lL
DKvFDwVSW+mDeuhJVqGPH7rAnm05Ox7s1ajfx9/T1jtBrHAsTpnE9z4powAro+oGk9LjyYiQeNbA
TeHrXqJotrpvyp/gTa+AY9X8KwfXOQviEtyv6i+UPVfTNYBjGn5AZi8soZzH/dEloEg63VAcHOOY
xJyHKSJeYyOjK80SxNR/kUOnO4z/rW2QPjulPveHci0d1YgNCfc7nNeCMMAl7lxGKSKOCJlghIvg
sKSHVq0KA3BRH0fVYm1kf9eROlqK6nUnOJYVoj3txdWfkcj71CFbG6h7Nd4pk1eXJkYp96uj7ar/
ZUAhDzfHRJFyqfiOY3WAn6ElWEDRh1wRgeK65jQjyXYFYJuhHt8kQ+SvrM2dERJZw7gipeYVN0n4
ARxOuY7+R2OE4XaPOZNxjxzhuAF5mUSMDordigWTPaqQE68F/SyIJAsUEG8t44ytKg88+wms20GD
6p3KxeSJ2k90hw4dSEoohI7c2RmwVyAmSvMLjY2kdpu05LipJfAFj8cd8Nsv/CTiGJGYjxljTyjm
DXbBD7qZFM9A+jeIaTS2XHwabnRIZ1VpcBZ8Jgk8W+WR/3jgd6YvyzdzOjl3X6+d6fub4hgV6flm
2j7Nybl2zFeVqUbGxeW5dDum4h/C3nB/G54fx8//q7TrXBcHLpTcLyS4wyeviXypqJdAPtssDdDh
8nntrhaXsYOQCa3zO2wVrZS4B45bn5NlIAIjJANX+9OxPcW6tRDzCNDLIwMsD02lPERRl97vCYxQ
fCaYqInzTTPsIg3h8/aSO/uxj2+dy88px8aoOfL9S8ORz7U8Srboqdu2RO7YRnh22iLQPWU53OOl
mOmvsiLRwRfnLeKA4bYXzUZCrgkGEmVeXhWb2QhUSKq9OvoJmlIM5A4Y4j1M/qnF7xEfReUsRMNT
+So7L5AZGuL/FzFdhFXoX5SlQSN/JeFuCtgUYuiXoo0W1U0N3qkoXXayPDfY1475OBDGO0jgQ2mo
rgvryCtjp/Wqs4niq76gFokwuUkgBEeivTXd0iHubGOgQipnjjXc1TfXedmBDk+eN5KDur7YM4NJ
/LbgOcTO4NsqAvRblmeJJHicRSJ3beqByRglY42Hy5ObNsxeQ82xs0n7gGQ1KGJXvXlds7u0J42/
9G+xcyf/cqETHAhXgR8MDlS6OJD2V6Ujig/CLsuBnMzyAzQVcA8NfJywN+JN9nuZ9eGTKh+9rFsa
EGhBQ7s31kOxbn0t7wzbsDBOoUoFxXvWYPSdtk8n4hY5ATWOkdjLBCaCOQxIvtLb+6h8oFejapy7
Ta21Ri5XTIOlEtZk2PjkUiXJithFQ+oILE7lKvlpBpx+BXW1AhzJU9P204hw2v8BeJQZmXL4aTbQ
SdsGQRogchfDtatTdxJFjKWJce6knunrf4o5VBAxgpAAHj0Xzf00wQU6eWg0MUdhTH4CJ56nYAc2
RuHTLJz0aolNZrgo+rnNK5hHkFKosVJPaAvmWB8Aewvz29QCMIxRtXGysrivY/o9dGo0c1nNv6nw
ZpIiCWDcXYdTiVFC9GCk1DYxQYB3cUuG6bfnGuGh55HVYv1tbvxTn6glKcF5UtbNqUalpPP9D+Q7
00rm+UyBoDA8m+6AWVjVwrUxs6u1/oVVW/IDjmPtc6rZ1c/7gOcidwAXBzAs+RURQA+1K81T6dT8
SC5oRKmEQxQ+Da08h2Pllfpa5kFBi/T4nzFxaAWZuh1Rp1Jq4IoF38UJ+7loKVniAnoq2f3INIQ0
Il4HnA7y5xlsYs4ooHfr7ja2rfjEATTk1LXPbQVOqjk1s2Gd7ImJfchzoJQSHbSdU3hIZxexDAdU
J85v5HVC0Ggw7Zkpb8owmolphE8V7MBBmcNiirLS3PvkX0y7UK4ChJpfDPpQvv0IF4uF5CKGbDgg
o1tOjQi3aV1evxR85u9BI1zhurvZfkaYzbhdNpY12hYNE6/p8jnIlQPeTssMNz91+y4ddVNydaW5
XH/+KXFujYSogC0hjN+gs8p8IyAHyXfq0q+wCjhNrNJRSOukJDFShf4RMw0sbTKCygq+A/zHRDlK
EW2IAS7jMDLqfKoXyMSHtfmKMDdvH4hG+BZJ3mc84W8mOTSSO343UwPvNygAu9fc8fOJbUBpH8w6
rpCTBMJbzjwQPDfThRxxcRjPB85txfficVIPlg/SBivVnUxw9DApyAVHhh5ae6CuRmnXbjojCNvK
NcWY/E8heSj0VGrLS9Vo4+VbuVn3ZYvkoyymb0cu+pwJJD505T+bA9yxDJHXT9Lb8+D4FO+uWu7d
xb4jKmNeXmMistBlQwFlzhaONxo7XpZYTJBmb0iKMAQhzExP+URUBOkAznLqBS16kLffDJD6wMrP
vVP1w06vmoH5R3GfQfIg0de+SeYyA/qMw5pJ4wKP/aleDFED1WAAOxW70IOGbbNUs8ekwRNq9T1N
5lXHC+kjsYpt24bVVdZ5Me6i4Ihwbdv5LzNX2eOlaIZUOz5KJV+FyQuUU4d9RJM6er+fLyorKjt5
CNaLUsQ2JWYf/llJSGrZlnx3eGsg5eiwHmQiZwpXr2hDUijiiBukuYFZQUBo/0OFbY317b1V4SZX
8fJhMtonjIJDPoRPjeEAFXXvlScNqdb5uOaJY5QmI5PGqbG8SpoPi4iOZmKDVs/1+fPh8YE62CpX
+iPYgwZpY7tUDAiGydRd0TTiY1m02H1Y+08IV66wVrfuRQ4bUqstaJF+gb60qg083JWqjJwWZdZ4
r1QJAB7zbacbVVRPRkUpY0O0eM8pgyELCwGnFh2d9JWN0QS5ms5Xx9YgM63Moi5GVnJ0Im5boeSz
PQCZMiYpE2dpzxnm0HqVdoHFBWJGLJMfwlR8n4e0QgesgGV4Dv+jQ4KpFf1cRB45PZcQEKxJfEHi
G0Pk+q9G4xVBB2HXXkJd8UFAW3LF608uv/nUMta6AbePbibkeeSKNOhIW6Er0KscpY9RiJII1aNj
UR2Qaqq3Prj0quIqwtFOp/jr6BM0Y30q88QAdPCTNGrlqsErsNNsr460KLec+4ShKbtETrELm5og
+Ti2Ayr3RE8aK7AzvWC+DMx+eObcHPJbltxJCNekAug+dpWAwMDlCnUFFAWBp0g8Ehpsc8w/nhoP
WI9I0eRx3hh2XznU+K9lDk/hbC4rYOqHg43JviiXsJ7Ve1JVZbpAPZJjvgIQe7bus3OON+Y1ZFxT
olOUecnGnfV0QJxUKQXP+7vsCZJsc6s1DHyWYQ8IyU7VkR47JxSGGMYzBmeD6IRqnhPzr5pdVLB8
zegTrs0G97hVN+EdAMTa1UOtM32H/3SjbjkCuZsZ87IvoaxQY27OGRozVIVQMZfFDrVm6qMmgYnj
CLtitvGzixFATbTfCx+t69V3FH2D8eLIeI2oH7y+tZAXgQBX+um71MA4SeGP4NUFphzVd4J2jRze
F13M0ew/iox9WrjnZnnOZGLN5M3xPDzI1OFzMj+3Ru7OEHgH3AkSX5TY+ItbTkNIbY0EhH5Sv3eT
Uhl5JC0iFwnBEKjucHu8gV/n5DrIVfyJ+TXh5mmeMJ0JLxPknVgHEdWdTEb0B/OB5xqhwRmLRnQu
30J1P6gHpwFbF0VpVcdFQLw/qt4K9UerwTtxhFiHMUbvfXfCi0UTD2BMc2gMWi9q/HaeRUG6mkcT
QmGxNj5Uu9ZijfCNwVr3B5p/EPBzGvQsTVJ2pMb0RNXbKFJp7+JhxLkLYlQTAE2gVCKOZkWLyINx
LfMzKY6UJEKJn+xEsfWQHXx1TUzq9Rh2413r48YcxGv39NTSNfGFLDnqoOLcZa49XMw0OedA6+9L
H/If9AthuAhEgO5pbssYtcupNnu90wZve82oe53yuLENTYvf81Eotrv1qSDPgOp3foMxj7A+IL9I
q7Fvbe7YXNx/KXRrS/LJuqszPkypFoPpEZmGUuk6rZYvqf+BOwENPRJ1b3nBDge0+UwcQ1NT1D0o
1XYV+H4bAho+IbPFGzyRDOIDpdlX6L3/sJ8E7+0120Tu8usex5VCIZ85/l9X53+OgQ5vX5X1DgmK
0neqELMiOkheBG3t1QIKec7YjB/XrgVywcfvVg69Fs2TRjYlO+towKU5peuqy1ejikhQYFJbHbJI
Oi2eqkcO1aVO9MTWJTWdaY/DExzTGwIzUjE2L2ob5on+gs/EOsgy51SgQRCY9VVPE1mql0DxMPG6
jDLly3e5i5Dg5bj7UPKKRnPn5QhwO0A3YHrzi+OTvc8wiqX731PNUqIRpO1ZFzCMNPkqsLUl4eRm
pXLQa7fqYfxwS/sBre2az5uvHR28zeOSnIZED7xaU2pP8zWz60HXj3Y0OESX/645xB3bWNcC1U4Y
IRbZx+gZGM6aJU6sygbHHQ73/qDApRYGljjWXMpSBM5QlYL2xDP7LaopGX9V0L6daFVU3MT2xlaI
SVO6GpY5tEWX2Sxj4sTCRiSN+O33Eln9+HZr5cDwqKKky2tGjbpIYE6AV65c6M0p5jBxgmFI1G+4
EfeS4kXLrcd+WKKjIxg9ZI/QxD9NQoq/cuX3MG7yRqPAoxnrtFZKsybQlgNCjL2xfJgKxXB4UwYW
B5kkCp/jS2OxWh8jJlSWgx2G7y2Ot11Unk21WEiMNnXVYl+rhXNcgP2/jaEl00Ea5xI19+ldHfkf
A+9RTMTkV+rMQopZyREdp4B5FZvukOd1sEY0q2knuSSv/mlx+pD7f24R0f7SBfPN1YjtzBYaczXS
vmjhLBoTyaagsktZQZQnbiD5wcF7OQCNLnp+cSQjANjp41Qb6DGTZBKsQ7I6pA4y9yD71PMmPoqP
zkfW9rm33u3JvwNFjJdCxQOHh42BCDmjJ4FoffF0DtRCGsBp0KiQjU7CZGPRT9Yi88WKcXKcrS+Y
CurLDFuvdOskOQOlfMoo1U69OW+xY7nroFAd45YI3+PeqnCv9ANLE5gyI2lUvi3UIv16wMs1Zbrd
jZP7bjMJWnwSmtdzfBxGE0uliSxwT24D2TtQKmdw3O/mcf7+8jwivLRLRiZMoZbMDShzTj06nYxX
ScfJuUCLV1fXJy/yQ1OkCJtNNftG+ZbMwoFkjKru8/61LH2VijlRc3/CPD/6b0hNxYPzKrKRhwJY
5g1lq9UT+v79CUppwoiBAcucredvRYoY1NztLYfgoVHB4qoHYmhfP0tnRuubDozgMMOmhmvdcBIs
+qhO7dk7cG0NxsqwIdNYCcfXe4K70whMjeUWqJVY3N70esLH+gRn4plC6Z5nEX0aHGB5JbTbww/A
5qyGDJ5zgnnc2KTybgvmFjviD8jUw4OHIreGaYpgSyV8qX51MfIJIzlJLQ0ByNwDy9SGClsuy3wy
NQNoJr5lqRnjwcKtPakfV/lQwHckTkrUjzXsxgyiWFa5GvfOeXJgipvO+5QI9lpNc/uInrLuio+8
n7vi7CTA01mzXN/Rf9tYi01NzJjJsSnKxD4LNVovYFEADc+WQyBf72R3773Z76kLzjUbC7TEfLYn
vciAUv8D+x/YcX4vuDhNbN/ZyjloDFHWcaJ9lWhDlq9AFNMvbAA5nGLj9lUYcG7uJYUA8CSaOmYp
ioRCiWXXjQZyZfL/6f/r+6/kNu3yp5hITaWPIGLMdydoKl/P83t9l8SOqBMiwDLXNGHWBwcGC9bl
EUY3bnrapXe9TBSuL19WOv+1y3/vkTxFb3QCamiTLlsZKFHN0oYYBMpsDDijGN0Avn6sPd7nmAZJ
03N5+CSo2OAJ6Rz77M8jcqQjHrtjb8rpQ301NcrILd9WKJH0iOuimGWISDsupkL8McXuHIGexFMv
aLcrzWMFbzocYuK5cxPURcR5ft6WH8EOs2BNpoL5/wBve3IoUNa4jssxbdoISsSNaDIcMnCWRXHJ
VsBFJ2DU0w2/Zn0e6n4Oc/OMJ2VUOqbpjFddz68pnSJHfrMfCjBMQYlGeZaEz05mMmj+x04Xl5gt
NumEXNsHrE0KrzWoe0DoYj51Lxia7ivHHiIS9KVNBJUpGXN1bjJOxkfuUuGjdw21lDT4+fPneEPV
S2k3OwjQyyre5mnP5MypTeCzyeMaj8IDAKbJ5O8Gm9jBbgO1VXf8iGgAm5CNisBTYkGbOzfRn5eb
/Dm+zzqO7COymOPjC+do0itcypJ+623joBdGXSdhr9P7gtA21UYZXICQPldzIOTQKVi1QM+8kJu6
mkg+VGdlpZbECbIE8qbcq+cZsCLoNiO0y6gjpRASPML67ZjOrwI0UP/1Vq1nSIqXM2h8o+ypEfNV
FTJMKwAMiomqVPiy7iR6HecBLJWw9xW95Sx2gKqWWzgkUV75nuO0zAOXi4po+rP1SW9fgzu0j4qj
ylpJwcUnZqgPE4jyrFgavHrE3ebr9WALy0Fc6He5WaDaOOwKFHnBI7zMsvezeFiGKeCpfoughn2u
+qO/1Wd412XBS3gSj3ZWP1nDPxzfTY7i7Gw5JDgJ+Bny+Ve7qa9G0lpbqd+AKwbaYgQEsoKUx3w/
s5mdujPLBFxVnS8QjR4CAkcOQPzeSdX5R5V8vWB49Reco3iMF+PrCMk0f0e3KdXsxyuDTmLZLKC9
9/NxyhOWM/PQ9ZpsMtQcqVqE1DnFhaDR5P67lJN/0uovER7ivyO8R+RHF3v+VCOiyyg3o1GH7EwC
ejQjv+K/gmW4mpoefx92met5jQrXF0240el7leKcYCaXsNtXfswyEebxd5BHtVhNUCWX+X4Ou9pr
to09MC975IuZCmHllLCB458w/vAhBDxWT6fx/1GqidpxqVBPf9rlIEIqP2nNH84TR6uxZfX4NOyc
qPfv4fwoZoDWQtgZrejgQs4Nhj5scXE3PLU6aZCKTEf8Ksbxkf4HlUVJgCe/zqJ/Z/QO90cP7tc/
m09n5NnwV05HtA07qjG5vBwqdjShFAcBBUWmN87XjZLKCpueTjQf9Gzzq5lsJB9ORD4/eANUk3PD
OVepgePsguEj5jb+L0HJq8vARwCNP5KRgzvAfl1cLzEQeIVfZyp3OOz+AwlpwZ/1PhcAMHYMSgNi
q3LTEXS37ypHabXb+ShDsi6WAAJ7geMv1OhQ/WZq3dB+BD4X5WNkbxlu3fq7dUao5WiCFwo2MImF
+VmB0a0OUiv3X50kqdhSJNTZ519wSQ9acFqGTCqRbn32VnAiyjdRM+wKDT87N+rQQ1heGC6aANMw
zjNeOKGKwDv/NAw4OBmwBilNBqKkQpg7qtwQ1EfmdmmWkoS3NStyr2vlHvCzH4U8xd/+SKRUAHHU
7HF2t7tqGPjEm1PcXEJV2E0SqGNzGQpEoXiUPqxB0MEHdsIpbbebjg6I0p//HeTh5ae2D6vBaZm3
PjP0MEIMio5wK1KazLEz6HN1Uka7YtN1VGb+NBE8Acg612JrrluSRGdp/W6ewPEdtslwlDcpTySX
MO29jALpOcKKn6gJaeGfP0C/T6l69QQ1BE6fii+iiBxjHGy7yLwwKfxSQM3YDQeu5ogzmo/JT9/e
o8ik7HbOpwYuto54mlPmq48DKs3AFBkPRB/o1E72mD6AH3Y1RBDSd1wwARfFc/oYYzjPShbBW0jO
mo87OBtY8qyday4M9hneRIdAX7yzPDtRDreXrykb+LmdJuhplpMw0Hdc9d4SnPTKeeHCg8Gxd5xF
z7Q1zQQhM94Dc98hvk1VWveCxcoYwdMVjTU3RDVR/4jqlGhYZMAl7OWo55OJo5Gy6csvogkBowfp
j2e3iiV1p+IWyVJ7pY79Vsn6tpU69nYvInRK7lBinHGJTBsZqzofXVSCJzW0VRJ0Z+5dagp+Ksow
m4Us3jWh3XUs0MSDmNzlZDRErTZssAGhOIB+bI4ba3ahRjT0az2cNPQgA792hVuXO0lfyci+lwbx
FYWh/m+PbegqN9NTfCCVASFMnlgtBmrXQAtPql7R0B0d0WBj2LqL/kSjkYfuBkN6fJ/ex2jJhgYN
dpQTlHwnXs9JPGuE2CNYBogd9Uu7sTW4ccFouTB0qQ21DZ5SOOH+8mWBj9OlWeIAL0zpiXjveD8j
qdQ7wwuLgyUKGAuAi4GW/WuOyFs7z3SHQRVFt8Iey3KFy6fCuk8DItkC26Cp00Bo7KtaVmL3TTej
m2eQFhF1ZTIbais9XCluQV3nVU6+gzMa8aNLS9mqTN8FKDJ5Gh70wCmbyB0LCQSj0s91O5Pi7Ri7
EcMZ4Jqy4Muc8HYU539cefYAQUlbYcRn095ZSu++DQoeCCywnmKKXEmB+apLVlaee4G+Q44yJGx5
bJX5uXz7xWJjcqzWos94kTAXCBabcJKUJKaotnzUAD8ITG3npr8sjVbwHrJgMYnKXwGFVh+Uwg6F
ETcH1LLBPPFiag+1ldfn5XXnufqwDaIwFXKVUZOphfANFEnqOr8ucuXaDRpylVJPj3qhWARZZGih
oE0CJcAYUovqK0va8yuie6vCbm72+nHrmwsCQ7hcZAHTr14iGMe7pM/cUXdo4vxV8p1RXg685jA7
IMrT08IFCy776IvlBq9La/umkIDussSYLZovIWgehdYU68vzTxyGcl04dnhOngGFPTJSDp2YN66R
EjK3W3mTja3CsYn8huz98BcdlU2HV7yGj74wpAX9VD/5e8Ri0QbaDdigZyD2pxFtwI6pVqrsg6mH
HPiFeAKKsmYWahek2jTEdjC9nw77WKCeBRkvaUfssQ0U/wx8lVEGmIR8z6WvdPV0VhxM4/Mu8O+y
DVyUlzavzhQo5NTbn5gjUHn2KyQ5MMKK9/7X/Ii32R/jTbAKCUuzWQWswBADMXQTO5xStY9Tlpc2
LmJXVsQxAn2hRtxIt20IYdvyHVuWb9CU+pqbJF+6gmlRx8byDz6Q8SyF2t1/wJDNfymFXq8qshH5
H/8wzVpBGpJaxb3Zv54QKRQhs3FRCR/e1SEAqmPmPbaaGC7D6bkyshcy1g/voYM+bvOu4QU84qAw
VQQXTae7UClVM0i3yG6Mu2pUYMoryU0HjWBoUesnNqUEk5sjLg1ic3N6blfzDoWH0v8Ji2U9oiDn
PLnGN9L+N9KU3EYgggbdXFTT5rukdvRLEFmMECljAMWcHqHxkt6VuqQYqtC2EpqX1gQW4F7l3Pzl
r0LdVEoTjhpUIKDzlpOu6vKoCdtkKX1oUcYbsiqt8TX90tPCbRlIKRWcNaDU/UmJ5hs2ihVb+u/+
aWDGYpn12p5wO7ZP/DGXmrPHVuyTTzoAvhYneRHgOUVvfE6YwDr13ZylYYAhYLEjfhw8bQQcya7T
DKSw+VAW1l5nobBLWG6M3NBjxb/dOoTQbMALP6eCkIS+0JxX43lUCC/99yi36+x2GhkSEswnd5bW
TmGanYV/SouTaK3EzB7OIETglPezt4tZcWYMHq9xzpSpfqh3Fnxh1pBvAQcjebWNpjg7NDuDaXEt
8W8MSfQxqvXT6DEIeQAFO7haM6adZ8hsUFCgY2HaXSFeclbkhwL0ZE3qdIPl3799v5SYVrzlhwiC
8waoUyzXVPNy9Ng3u1vfUKUV1taMaV4SVT2G9d5jBeRuCEi6GTdAh/Zv4MKBxeImpWJqZf63AAtE
SVu0No3ZQlaouQp8NA4HHpLz+wXc9sfA+NgLf6vGIPbKCuHsrKr46a5GEvDOkVWiXLoA+aCtV8QI
pwQFrhqDa79rLq6rwX5Kd3xxupsF8GMC0h6eXn3Xjth6yQ/c/qKyup4VQ5eFDamsDMRfQwtMMSCw
nPUUJfAMgZywH6MDjc9GSNQseIceKLt27a5Jj0D3BPCFa9xmygs93Awnj2oUPBNKvU0/jFXmGXbp
2AfLSeJLd+dhvBOvfmRnYP9vk/ZA9ALJSGXxlwS7YAHhypULJl1g85kL9E46R8AcKYzN20jUvwCl
m6+Pr2G1ED6QrVJfaoUFE/97kfTWY0KgP8PDV0d1jdYNe/YPX6lkATy90xUpIFqiNsK7EF8ZWePW
JWvOpu1cUVyFqThWjWgorS1n3GOA4B4ey5UYtnUKButmDlVWvImuZ6Sdahx67fJ/1bkrPU9OVRym
VPoxDB/EY0Yb34ImizPhQjzMv+mSl7wZ6ubUkqN5MKtbHayg5SiQQFe1fbvlB3CFTiuYO444WdO1
zCYKe/vDEx5NsoXjHvclwJwyGWlpxVMd90zrjBJmT9DYyU+PNvCa1xW5dxF3wIMbSoRRGeeeQ6Zz
9cM3vNqpSTFOFJCAyFqqQrjkKMcVvuI03+4502aXcLkrc8mpQKLrlw0scp1R8QlDlgsaaf1E9Ze9
t/hlOEULGWpWIvtR7Yu0Z+VierlHD00gSbbHKxJfZ0WwrdblmPVNr3SkXVcuIkzWvZ2kofmdepc3
U35rzv/JK0sBsDVF5gFBQI6HAt6Lu8HWwVr3eG9mdEyjjhr3700dWrTg3Hsr/f55ZD74kINCnLAS
IHu/J2LB9ykC6Bt+u2DtM3iBPPdlpX2b3rtt10fSq5Rmw7hLhcS3AzU/D5DNksjEjSqxQ6PgHqfm
fguff7ogcuR8XeD8FIplBqCf4nEgs7sIzvR+PJrxer38jlH7I1yYaaWPqXX2Ax7aMEGz9H9Js6Ag
jBSj2CJcvp68e07HNs0GfkSSNC1I3Eb6g4r2STlDtMPCqIqf+A19uvFQnRz4fwO9bj61/0e8DZ5a
q92Gfd/zQlHe6nSrcQrjmmcM5cZ61Ubt820oCI163t/uKnjJ5HnlUXNpoXERTQQFrxVhGhkNU8Pw
SlH+mtlXX9WJarBhmHSjdW3OlroYDV3Lao4cjZJ7BdoL0JKD0U2heeRA+PQ9FeVzxO2TSsFxJslJ
bFTyMabVMRX8NFeRefrwQWEcTN0OeQroRgVB9KgRkyqh5oG4K8ZENx11V9f1ac2843zN6mzaw5w/
5ZVh736DmMv+o6Xs5rAuqHdsX3B9XFDFrVvm9Rxa6yLDANfox6n1z9rezTrSgkLHIyzqN/wvMlPC
cnp1D618lgT0U+k8rZedA4kn57thKTP+WnoEUfeZxhAnwyMSTU86nQ8aRfGB9kkEoPEVGLpgwGlC
6yD6xXUTk6SNA9UqlEmuai0KaspF6DocF5UEtFNpbOYBITJY6NAWnWtYEEeBBv5vny8n2fmN0i+k
jCMypotT2NrVPOqUsRABmo/1kg6X/74cLp6bQDkbqnsJF7bW3Ilo+1S8j9Q0RLcrgcpbXGZNnyWz
gUawMB0pgvgSkTTsQ8AfvskaKMQfGPeC3LhkWL1MNnYIFZMEyE3Wj+dCYECzDSU19PeaHiGk5Eoj
LvNSBlTiZYsWiQpLHL2vRCGNXuqiYmOvHnQSKxyPZIaLe3Vz3klgUzRLGsKzazs9W4xnSN6uXorB
JS13CAcnV43ZYmHDHtXSSV9Lgz/3W4QbgqDcmWCbG/q+aEx3y6J/txPOgzzkHL+keNSx5zYhsS6/
HT4SRzJOlEdmw8iXYVxvZZVm6SW5qJG1bx7pH3h1weI0/Eh4LYsrtc48r7RtsMtHW68G/F6NED1D
bwt0A20CTa1G/dyXT9/xp+ZwmmjWWdwAMnOcOfTjnENmYOFLOupjV8yWu+azF2XeAffVpe4IxOBq
TnJ5SL/6KoqdW6oqILX6+8BzPSo/FHKgT+gYn+RE9SvVaIYotCKdV/UMIBmxeRxFtvdut+xV+WX6
6U3BooYKGE9xkxTcMXM8LGYrHksv9UN1gOG6YLWQVwWKKfR2t6+r4NaQhapjEYfXsMD+st4gI6iC
7ywjyj6SgZzIfK9tSWUId2omWwHvrf6AZesyxqB5M2MjbMhrBZV73rxhwJHENubAjvYxq6oGP/VP
BHhP1oZMQTaW7Eu/dy+VWoWtof3uNR6MdDC3tLrhsHgXPzJmBhxL23BRcAFtRvMvswrlGTtiLAGJ
K7vy3uZ2wLoNcuebjP4HLRROPdpMVTCX7K3mjXBrOdiflS70B2tPqjJcYse33fCJ4Bhdz0adq7d7
rWgUBAyc0ueJ0fmA9V3UJIuv0hbc8Vb75Yi7KZYsAe+jUbnfR8FXIpUAbkiMaue2rd2H9zYD4qFK
XBHI8odngwQc4eLGgQZhFzBCQkuk28oq0i4h75+AyvPxsNs/1wLukTVLgq9gTgxMgnO1kvVyrKlZ
IHb9iHpAZnyco2CgqG3/s6MM6scOXuMCnQEbvYpBy5JXHdmyhgoXngHBKjAh3P0Dh2DxYm+NRLut
zfdAbZih5VUydM53zFPGaWwmGlabf7KiDpNohy2tjLtkGoLLVUQGcezzWAOGcNCFe+0LJhLipxnY
gfiCJcfy6TvKe3fIEOMq7vKeiDUrSi2Pw6cdQRaToTLAJTjqr32/k/i7duDOaEH8eFlveg5awoGg
jAx0oGdrvSZJN9H0lpY79JSnVZEXx46p3AzyfzhSN3m0C6SYWDqPMkHU8r4Wk3v7+hjqzXTa+qof
UuCijReAoOynTJNnkitzng6qzRie3nlloc2huhhcra00Fmus58pi1I569owT+6tqaUwLC08xzizq
cNQ/YLjNq8S6lLT+7rXCwrxkqd7tEhSjfMB2xBgMtKII1IiF5Jwpem8aLJN+4ilgkYTOo5xGKyAw
bBgKOHzV5ZvrLyWrdHfIaUodEqskzSWIQAp5PWISJ3yQOsZsPmX3buecik5Xe3vyepZ3l82tg7k7
k2z4BI8voo2pNQJn4dtZpQ7i2+JzVMBzl9kPDH9S1bgdEf0xEXSf2yxFYI3omq6rSBXc6I9HOYxT
0atgasiNj86FpR+aokTpfdPMJ4KnRlf4STXsXcI0/SOs85ZDDW5dO6+ipBzHh4LKdfRuJrW0dtnt
7b02MvJcA+SSiuIV1S4QfSa5Z2HzBlp3j4B3+pEtTVzlaolbgrg7oFQvjgkj4+VL/zNBWCA96YZO
44crj6/BqsEXq2QEJ7QfBw1FeI9JUVdsgJSPhOkQlaNAjNc3rdtbA3rljpXnBvqhLxTGp+zKys1e
/EzTlc02XJx3iIQGu3+Pn+Ae/PhTFPPfUMIk/KvwcL8tHiU+EuH2djjxC0GTaAX0DlIcx79tPNwv
041gGCjQW1FJAvnKKKk++0mr5nX7AnzmHQDjBUwvtUNGoYUuEE89X1yOo46KinBMNPWdlbFEGLQJ
cBqacfQOHzr+XYr27uL7o3XcwLPc+uzWjkHS5O/aVpC+lrll6/BCxUJiJSjcrk5aFqKubrjpigYX
alzHjJQqEeg/ZNAg3JOoSxPHg55uJjYFR33I4GS3x0FlNmP5UXV+arN8AJuAm8iOm8Ak295XlD/P
Fhlt9wLrMMBJVMeYrUfK8wr2IL/LQhw5VeE5j4Am4ZaA9he5R2pGY2jBMigOajlxicEBOdymCJkk
ohrbjU1kWS9gneogBmnCWJknGRx585/ed35hI/rlExWgGjxeWM7pgBACBIQGM1K19VozpJzJKb76
Wv3Qo8FvjKe0ZF2zhVfeEtiJ/CcLkqZmbbUWo5i1RJ7prWU8ExX6gUPx8Tk6u7FDwWQtppR4JS6Q
qxnwC/9rFpsHvMOrzuaCsdbJkd6F7k+xIUY7fytzY4ZPW+ghFgb0rB8kYY9Owg3vjp4HnX5kicCL
RSLXuIe3C1/6W2NQyBgVMPNuD3oMdzmYCWTdNHG+WjS0H7MmN/WoXj2oVyOaDTvtBzvaA74Z7OFC
PDL9uP1lonRJ7gaPjOS8hNDIpyWSY2KpDC8Oxfm3D9nD0+dJjPK7ADqFE6vuE5a0MY3JfdQArNDc
cTzTtmQc2RZ9EzBMwLo1unG0Ql+VKL6S8t5PIGCDZcbol09p3YR5tAWQWi8heGmPw1Y5VbZn0I+6
FUEEVHuUE73gorEGEpAC0LG8qXottwAIy0J99EpHnLRyTSJANmiWIJtsfeeacnoSN6pqviaQh1mT
IO5y4WqPlPP5XThjCEqRZ43rR7bRx/NqC7i35QGTDoIfIUPoflq72v1eX3gHD5E61ZKKrOAuUYNb
sO2tKE9Amb5K2Biadf0/mzRnXZ4+NUTNnYp6ZHNS/BGmTG9wwBSLQT+gKbCeWW2AFcVK1Wyy5Fxd
a9RrZMjo1KDVDq9vIyQ+4bPnjRllotv+mrMSfdztxGSXK6iEwdSQSlnd117sl+CQlQ9jaDLLz8KY
A8hJQIXr5JIknyqQDnUFukFzwTdOa22wnuLunU/mE8cKqvavX1iMFUlNaWi10mYsQJGXUeoaqMBe
+/4PFoBEjYc6yl419gpJO5IigfoMrKzFTwZknvDR//H1FN56/KSgbyf5S71S6YIb62AV032rUdjP
tqLZlB7SFomwqT4G37fpz9s4/vKTms7HL7elz9EWkkUEgAFjAhuGe+5fInrmeWlo/JU3390B1gDx
H2URefKv77h9pxuMoFTPmzVgPiZRUCT4FPkc5L6zFKs+G8WgC49/+k+jefvTzXbIcdkwJiPSopbN
grEUfp4AXeErARYQ3/Bm8Fgmkqvv/gb6kYuFgx+sGnMqGoJBrIaNOMC7KN50tD/RO0UpGiZcRur9
sp9kI7kzSvTDTQ38cr/l05Q7NnrrwyKXwqGxmRYQb8sJWWUmBw8I2IUymXHpMMd6uTwW00Z8Mr/z
dlMcMKoDurhjtPWi7CQvyYbEZtoKf0sbNC3oXgDFBzU5XEjmfQ2tOQyQAW9pN/B4YlCM+P+c/X73
xhB1Iofa5PEXJ4EJO2sn5oDXS9C9iO06Lx7T4gVXgMJbWb5lEFy01305DsQyHQlji/VcZ0cobaUp
7lZ4jscHHQwCfgAOnikzMLUeuHBZsHv/2h5XNwmvQVcoXbkRtsviLe8S6q3OAdksjyqbn/zndS0D
F4XAHDybljpNWZAceRrirWJtt6+UeoFwZqFD91Cv1flaVlqTMCicDgTCE0ikm8244+WYFeRT43H/
RiHhWBucFM53Ml8Jw3xuYra8ChRc6LyhgqVs8a9gRbAhudGXLn6IVUNPze2ItmwcIW1oEGCqSP+k
t8BkJHVaNFnq4iCzkzfB9uy3AJ/Es3uCViaM2SBkUJ3UZAb4S9INFN1z7tiqH57dbCR6omvsA7nE
l0q59li8Y37MfekX+kHfxamlVln10giyeOciHiyAh2n+ps+Ep0Ec3c++6C92hSHEqyN+I4ycddzX
QKpzU8orW60VjPgTZNpTpR6j1GuEAiUpN+P07ojgpTSr3rCHT378MYPqHZcD8VY3f+78x53Jqg26
KGDpoqQAGLJ2yXgWwhpB/WRNvJPETPw8MaIaBCdmgSrnVT2F0CNoXE67Ds5khkBcTAxhXMvHiyej
X/y9DLnZ3FGPIusUwWbNyrhnR2zjiSpQvf+iU+kPEt95qXdbKXvpEW6M36WFU7oBhFsTwiF56Inh
hheAWe5In3ybZdxHvMrb7mTWo8YfxuaGU9F89PDMiD94xqA96F675LAg5usPg0IIKCQpH6iTR3p7
Yt18gYdnE25Pm4ZAXPyzogcdCjeAAIq5i737OdRolttYwmeV7yrhjYo6yaUMW3YKC/MpndUn2lw+
Ud+5sKQ9Q3ftSJwMElWKGE0HA9AsPux5WfQXMtQ2ffkvQP7rMTihzP/F2L67PVn5mBQe61zRMxyg
FCUJOjNn9SgUtIERDA8vQ6RwpeUEyZ7cS3JuPv25Or/9YExSwDc8OpC6E9h8p+6/hd14h4B3L7eX
/iOiO8P2q9SbQivzCRsEI3zHm3QZBP1lWdmnfU5EZKEx/wd85fPX+j64y9m/gcKheH6Hyb8D8Jph
U+pOiKQlTy2QKLvJlwUzVOzER2bXHlWgVvZI+/I4j5FZLDLa2xN2hZedkrWaz2hW5L4woKTxBnIv
TY6iSYwpRSU4Os0flV2UODYzLMZVkkqvsGfQq0tF1xc/2Dir9HA8H2zM8C7cogXQoRZahwlWpxAj
WgPt27V7K1K7wYGJHOBAU8SdmWrDdUNbNGn+cOgzdWIJGzOfmHsw0O3xkHa+BCeuk7VlqrW5wye6
mIOdN4RrrISV/Ivl00kHgOBkFdYFln6qvbD0C1WyTTF6V05qFcwJ3VGgGpYDFpM16lH3k+P6SM9v
7yCRFEmXt/q3xD2KgZASefbrRimvDL8zVb2EGN98k5dQBBX9jSUsqVJnrl4VLeb2l8+MkTOh3L8U
G+EyKNJkTN+mIgCUPPMNEDkJNKPCjLt+IsoUYRnANmAKq/hb9NOqW3rCFd8FSM1Ao+WV/lbL78qI
hc+uT/4QcrtRTGbkdmednw2j4eTpj+Ia6UepN+MYqJetPs/3je+Mu/938mQ4aV61e7iAOuwKlFMH
JMyDTOwvChUzbAJ//aa63BWbCLnNJz6OeedVyncnm0ON9w8PTiBUek28u/qrP+fkZoRgUWwjLzMM
QAgZvSH3nzcJZQOAyCu5lDzksj0i3ym41JrhfA1sRRETdFrhr6GJJvA8OvNppccMOUYuvdsyo5/X
dd9tmINHQ84km2IZCgtrSI9IJUrIMczlCJHtyS2wWERsKX/Uf0icCkKT9pGvjEo0Hahepzu4W5Oe
1CewtlzuP3gv7tkPr4GXmxULDsO+AQdLXxE1q+i1bQoWStMN9zukKXhtZHoCjn+89uBQNztt8TKk
l+NSXb2Rerv6aZa3XZOzsICSNO+L8gLcTmonkavq1aWm/G5xito+NASEJgoWaePK2WgezL1zdofq
cnYqhTUkEeIGMQyRSuMORyjNnjHR7pGsV2Q13VcCGJfcgmnXrPh0XrN2yRdpWQwabt8dBgLHS333
eMqoLE2XkyFknMm3CCvK8bAMinlGkFmBaIqV77m4jUDfT/1kB1MMQU/OjKgOnotzN5m5IWwiyiQP
gLYSK9IwqJPLBBRcmU5qzLHlpz/MjRbQzFnbzhCP54UQ14UBMp7Atw2xvpiDXZ1OgWU81JKZMg8X
IoA7yNdjY8xip7Z/kRLkk5LbT6EV5K++7k5mvd9+9VcoiAzWN8GcVHXh/w4+NNLJHhYKYAdOYL1V
zbPFbEgVyGkIVgyyJNg2Bh4lQvqoXkR1zBuyMRQA2ly0OAzbauUH7ZqWua3pDT+7C6gXI9lzmQm+
E7nksFL9j7RieglWBlA4RrZnJaWLunlIl7PFKjb1jklKPa9/+fQrZIgA5K1HImlCHxnEkCqtZ38J
nskQk2TsfljkTV/ZX2JKK6k6HggEC/yy+Vp+jSTyrc2AkWUdGAlnVuLHM8xnku39ihOVWKjZ7Uz6
x8lQBsGB6Tt/Tu2q8ITCYvHjT55nCL5/NWzHr27J79ciLuhNK1j85Hqf28R1QopBdHA5rgZswGIl
qJxer+r2TzXdJooEdtOwx9d8Gy/zSrGF76/4ta9LmdEE3e0Fp4aUCX6wa/5uMleF0Ytv8piEOhU/
B8UmYeyTJ6Owz0edwrcrFM33XJpGu8cWxi9ocoYe3pVaRI9FIJGVfvAteDZ3By/nRFckWaeuY2gB
BDf1ZjP/uroWnrRcQ/4QlBOiPTyvkIfKMTvs62z0n0Ahn77kkzNeeyT2GhOdtH7FVLHBy6mjxkLP
TnR4nkvm8PvF9hMNBub9XkdklsadriMG2fkzXmbRfvgKGzXyZA1ALAAChJhMXzwO9Fa6ZYnZPs82
iedK0n2nzIsxeMybCmprz5aejh8dRk4FzMZ/A8TQLrJ59WuGsKLttySTpmmRhKpDW9pLibgNboGN
rZpadM/6TS1tESSqRbIQ3iRdNptJrYimYv7CMZYkUh9KIbnCmOUHvjlXX9LynPxBrGlq/RJGwclH
fPrYjpUZbTXk/OBmxqElX3R5Dr+eGXTNJZa7U943Y/GPCQs3sOWZNzOIVPepQzubUyeSNKZ3gPeM
dVooRrdxmgub4xc5gTkfKom5d0W3KYNML2vAy4srngHJ+HkjgJ0Lxb+JZFmOYafSk/uALxSNP5fv
4hXKAZY4Nmx+GE4PnSV9EPJx+7B+RhsfkbqvOSNgt5d7zEjN/wjJ2DIfV20k2VATpFzRhSqzVfKi
c8B2qfCBFXd8Fcgvg1OO8wm3Y+B6IwvXfFeqmSCkbSt16moIb2qbupzYIeEGl5KQaGVzvt1rBmc0
fIu+iTb4AMyxY8yxqjAVvh4M6rkKzfb2xC27Dn+0vAdDOdQPQ/w0FbAL7kpEbZeleAenkCjTEYEA
Rh3JOpoqYKj9bxddWKDVQgyiiIk/AvKBsY4B/sRvBq8r2pLkfIU/sE43xi6m72jlx6SNLYIQjJLQ
kAf7zxMn1OOt4N5nwJPbAtmc+sIL8jnnzvtUyoyvy4EZG2BV74QwcnAFZUfHi5YPc4/z6IMRrZ3q
lCLVI5HiDU7Lst5vS52JnhbhkjgCp9pfg0BYrWAaQW46OZyVlS3SmdSwsX5Wv3rlQjmYeKW62kBR
9gUzNeWsTJ7o8h6MAABFpUQUUWDcLNz2fZNDL9lyHxjhTqTFgUtRNlhwCdF/P6JFhxEth4rXPKjk
++xwjrMhL6Yt9S8Kw3dRLk+YA2mRIByq8AueJyfzQUN4l9FKJX/KlKbl6e9Ds+ch0uV1FSAluwoT
7WcBdJwd3ZNUtjirLLaFyRlhSdaRzz7Fwsw87SE3F4/IfJOqmwyeLM8B5WSvK6eASXkz6+tAMZgJ
yqg6fyqrU5BfqyaWvEk6AHFBGx/7s4oJ5IRS/zAOyRUicQq15DmzDe1nlVHJPpFwQaNuUu/BJEWP
lfFEZv/DfnfWF1jIeaV8WWn2JSIopbOBDvYeqgA8TwZEXBE71DA52bs/5Fw/jsfcLFuJj39MOA4s
SZVlUL1eDbl3qIr5P0ewddbHSGalMfmi4COHok/gO+98heyzwwZ/3uHRbpzOFtQuYt1/6cyBIAxu
QepNAocrLZ5+DcyAf3dUJqu9/IlXJmYoWKMVBTEwLutqukBy4XxjR/w4eHEOqe+ihqieaPaWi3y3
qFF+5wZ/GqOQK4pFZ77uJjdm9qO+Nr/+cQPS1lWK+4C+iISWmNpqftqHgBywl343V1KUOk+/wiNn
CiBJK3swJ9x7S/nnTcqdQMH+VCKBLy+xvUj2Eld4ycLJVIIAzchoE/nPvUDp2+KUan42FUctO3Ig
q+/Kq7Tdg/6cPu3vO8MXmHqzx0vef9Q+Isd7REBwVgqfF1jheB4jqN1gpl3Lt7+hZTreFURxOv8C
3U4RioIDvn5pern5NH3HsMS0W1lbMsI5xc2hW3KOdk9XYLDmJ7tLbBqUUl455eikCep/OPqMesfV
oAyE0p3EA2g0ioSxZ+S/I47INgsZQjbksFa0LwNJavj1Dw66hKuWAaSg/yXu5QqjMsVn6WBaIgqp
w1EAf5rHOjTX3WU50QCSt0oRBozo/ljtSEu44AyRL5+J81eCkvYXJYkLB2vUpuBDMpuXphEfWkWJ
9GsDHEc87LSiDNFcdknfDpBg/8U9hiuQeUU4tMtuD9cRZHCxwTO/GOX3pwOZywEj6W9ezn0U9YeQ
NrCxZab1ucKS3mkPde9abb4zmWMubEu/kVKTzpN+KlH7E8U1lZE4ZrkAjs99WuUK5fNwhc4LWVo8
wWabCERsBjlPDjLKfZs3lV+LJ66TVBVa9mDG2xfU6iK8COkk4ctj9W7sq1kOWgBtb72rMVxaO9QK
J73KsgqQZF+y5HBp58QiWGEJIc3NPuioAMGG54eLXEreLh9ub4YhLo4W8fYU5svAtNmH9xJ8xrAG
4P9Nc4d2ImvCDxuWPnj3+PP5av63/VTjlVowpcPMaZxwEl2TGG6r05QVJL5h0i1ECM3+kjNs/Dj/
T8a5PaQGQ9reGanmWRBeg18pjvbAvBI4ZvSiiZWuqsf+0y0GjBZA9aHKkJi41gYbeBq5XUgKsJ18
CLgBVMopDgWLof2699o1l9t+fDr3co4XPO1ktN5yN3fgwSKVgnxtBtcup9z1PsI+tHzK15wBhvEs
eqIcO0v5DwGDFFg3X0j+Zv8bVmXOOk5ZeI1GeBmyQljPJk4OvwduWi4Kl9119kav/l4uISGoQNuz
UIk1pH98NeH0Y/sVFNr4Kk01ztq7R3k5OcmbetkRmuCguzNrTvws7lhtLxWpkc09JVYpica1nnqx
Yml50EKmWV9kRBjtLdtaah58qH4tcTaOtXxY1tlhx1HpgVR4K0AXNOQg3c+YjOZauWIUpnRZXibg
80bVtx5+GxBOp2S0PGpzn3xJr35dh0ZgVxuLnW2QjtGB+f0EbTBdJ3V9QcEiaa8DiXSMpyDO3Q4E
COEiL5twMqbe5t44TCCf5KxWrdifyXcYWwAXAY6Csaq3gx3xOMjj+woUzxH39nRb+Vv8E/G9JIh9
cbK1JixWUdtMErL/HM/xpDulFjlu/g4yjQk0wd76p/OfPlVHi8lMfSA0KHDFFQH3Gc5VjYjFZjGd
c+F/4bZyfBcELxDHZQveYuTfyKu0j+0knbU5lQq51MlNTmW5nh1rXZsBPtoeOc8x1HL+leU+vFiH
oMbhTkc1VQSZ65dd2X5/EDaWLIBBdZ0KMDyc4tdkm7is0xSlU8oVxYRa9LIrXgd8gBw/s92Qb2a8
5Qhlnu14+LbBABolsPV7o253t2A6JPxH6mw+pi/ZsNdf+e1vOIkke8X/omepoCVGxSAcAQXwmGXY
t4ln+4amqA23iW4gdzW3OCf5ijdQD5fG0j2z16aEN+0KZ71hEVrn/pBkkLKTaEX4EXPuWbO+XdLL
tYUgKsuauUe5YF0TXoguzNyhZIK8HGtJhrfpw30YpyBp8voSReu9hDcFeO9P5cm4rP1afiPD/oRz
MhVZy/P9rCwQcmVQCUZIY6V4UVEupxw7n8KEfbDQSYFcpjWm24QoxNneJh7aYMnromyRmerWWOyq
5pXczHynnQ+9LxxL9YrB3gjlR8da5BaG0OrmnoXlS+F/OCIzi+9IZlZrsIV8Rw37Ky+0N+F/IS0b
mkvRDL1UOtg8ZJzoen9KXFWX28az8DgrET67IfS+jy4Pehld5iNjAJ3xnz5slv5m9h+TKdBqLDex
Vq8oM2htCkec6MkGcWWUqK9UN0+r73XbQitEzgdU0apfhbZvLBK+f8XMCda3dPuqv/jbu0hnsiWI
V2Qr5E1/BXCxqwhyVsxQRYTNNBkQLwpNkgZHKym4fQE9RvvhHx+RLxRGvMPKe56DgcWWPsUTarL7
8S+JzhUi3OgcSUmazPbb2/CIFZICGBa81eDT5j8aJreu+D99oHnOMfJlTEbBvUZelEf7WHQm3q11
9vs1zvBUWKixewK+YYt6o+V7WJh/07XyJKBFncyCnBgwsSiwoawdnEEa8ncS7UgTm5wEV5Q1ZM6+
cui8W7cF5I6j/DDFNXHElug4ifkXBAu3uPjySLm8pWJUUHXbjlaBwvp3e09e4mdHyTMLxL950vsE
bfw/YcGzUvITC4tBsL/Is4kqCpUl8WfNFHrNNSoys6Zw0NVuY6MA70gae8spGPQ6h4eZzTB+9pND
2Vi74wZ2PFtblYuRp6/IyRwvM5NmeDCsTr+4at5uzGquxilt3VQyVuRdJvoBcxzZKS1Z2RXTjcKq
gppYbAkXHQh0EAilipxlZdy9AXBEAigTQqwehO3KSpdcjqwZ29g+mVWBkankqudB0X90YPY9MJq3
z/GmruV76mftoA8G3/qq2cCS6UP4Mva6KR3I3FSzGO3JpHoD5cw7Od/p8PojpPnLvcVK3fFjt4eU
uviRgNUkcKgSKOXoAQ2NyComs9jEHWH0kzikWdtzQzYazxKl4TwirLnoZhoohcGegiSoWeY1y3la
hVMvuQigFmbNkIhWp5KndusEAI3tz98n2Km1Uc2yIYPj7M9Tk+lt9dPc4kIReMqNp3ScSSWeI2xE
PXDFf1yl3h17DRDzrXK6RjURch2qZpwaxtpCEEq6XzzOaW8lq1VA3FmRo943Q9Rx2pcDTTq2LThF
OlXW8sEUKjZAD6vuBunt0XTRVueu3Yi43/teuws2YeBU/yT//iGV53guJUYIs6wWim0z2s5zFCn6
e2XuApNB93//54ymPWr22152Dlw6KIxRBUgZXF4xDYD52o0hXgMl+byrsOCb25DoPaoSVX3ONuMe
BkN07oYphsYkJgT0+v2M3P9jvGq9E8iih5ziXH7RCQjG8f8sDhhWkU3fD8ht2ueNgAtsCVKnLk/6
NxlM8zpByFzXHypmrRPZmXNg9WRSMbi9rkwu9LzBxXbvUjsmRNgyqCwpOzbgp2n3RitB9+wvlphI
d2AOxTt82gMgl0P9xT689VtAJ3aRONypK3Yjm+qypQfpSq9x9+6wFolqEHjxPBGPmi67W83ueVVg
SfcgZjd+vgoJgzi0GguUkzhihxFj3upaECW7YHjSxx7B0WFHI7zYVWA3yaBLAGMHBwOoOzXzCWUZ
0VUbaulF721zL+3++Kr276gdRvJzdLzFtnfWzpnM6Y1JGlJAjcI8nKvt/ZKoxWle0Gui7CxF2hVZ
bNGx05q2IyQ/H2ns0Ov6x+CM2Xhe+BRGy+dZIcl7h7zW7QIbAZKeoZEstsELQi63k0W3LJ0I3MA1
bHiODgXk1n5Bo5bWQ4dxBmdFsGo/zS7A4eDfyASQqSDmnt4RW+xvDZuYRIt6LMiDtLmX2EI2VjKD
O1IZ1Bo96e46yDPShtdSUrENE5aRmG4OfqEB+tiMDNsV2Jb2Xrn0bVPhyoPzu5SE4t0eQkJbJF2b
8otEWpdTK9dALXclWroU9s9S53DTkv713ZhakDW4y0uBJE1LTmhP5o8qGPHwS9njsRRgw7baDbkf
dv6NRm4vvpSSdczBSdxPbJz4xEnfvKz6tvx14SJEokkJcAzFp+uDtUL5TnN0f6xGF4CLEa4Mfuia
MJO3mCQ+c2JuFd5qCKOiJXn1pVJgwId7mmZEz6j4vaA83AV9e3mUwYixP7plmRiOMIA/IdRf8bzD
MTutnKPqX4j2ie6BaJ6dWkW0H+qyXU7zzTLCJf0Lis2qBVkwKZE9ADxwQ2rjg2LVNgOErJPCuGYq
Nhq/L69miTzxAdB1ydX/wJ/X3F8vvoDfauHrLtEvgHbMONhKT0EgO2tHMHNKlIcqSrRaWc0GXpQp
8zGoNcZ3GF6j9kUCmDXqbyqx11aHe8T9ZQ2s+CLCggvCmK5uP8wWLxZD207p75yUbx0WGeFf9oW3
qfvFV4Dz8wG0dB0dwyidUHxp4eFkSkXAnUBB0/bo9y6PjgPO6+Z/HlJ6diUF4CZA7daHWezE2oRZ
xQLkeOBWZ7nY+je1gvVQTQhwYJak1MXQLq+mZqXRUYMuvSrnNDQQHofV53TkZ6rZXgaFNlc0Ma/s
KZtpMYQStvgJSbAZBWYipfFZAq1+G89XaLLCSJdjELoFBq6UN0w37sXHsAYhrbGOqu/Mg0gc0ieg
Wv1+a83Xu2IRaIuqqYym77o/Qx4WszHl7Fhs6LjHcPJCfJUp3qb5BhscmyWRV1yn0ARJPcqAa8YY
TKmQgO4GKGmxqMA4bdzXpDJfwcHZKufTcgASpcpAuBVZRurb43IU5Af3DVagDB66zeIkKeaBBYc1
iwAZyfrcY9gYGxRgQ8f43RpuGQUjI1H1Xm064yOBB8Z6paRu3Y3lSmOqd5BuiEB0kcA/eIc5Y9ay
96eBOBz8MlduJ/yMl/7msGKVMsCEq5Nu5EQQG5zKTNs7TBdL0wgot49g7mbzipuM0RrmRj7GSkGI
A10ABegk6G5bmmmkAe8JkqdwT4MvJz+yXfcXqcKd/hb0Wtyj4aDtv3fBjyeTc2AaGSqQ6gkt0JIN
FcvuH5KF1N09LpDhcLnfoFIXzXJTLuTJr1Z6VxHqwsJzCvKw+a41H5KklEgUQ7BfsltRkugrykFL
VLFOC8IXpSb3HACQOqak12gETRnt7u2nBszEILoskDh1/U1xMDnA6Spd/N++ERBpnXhPhXAmn8y/
r18VmhbrfY+Kq+Twzte4kaNiry2EK34SLDBK1YCm039TIPyGKETNTuEHQn+ejebt0LbWv9GkbAJU
50CB83YsrhpicbLOmxEInoVAmkqeCoOJlCArJsq43XbOd9Z+BQ/iTiAg+HuXCl+8cV6LHrxscuN7
qnKPMX3l3KraEBYS2o9vceZJhF8XMob5NRxr0Ws6plbWyySyczaIdOWX24R9GcPuLRkBlTvePgrO
9TcVLzlifVhIxwX+ELacwkGpq/RIbPQmLOnxWVHZaeI5ksB7/Wj1Dmq4c5T5OQQJKfDElGpYHDTh
rhciaOCWLNjWoq5G18QUa1HYE9rkkwjHyyl+RelSBi6JWiEveksX1jM+1PkfHmPUq7jZmmWIx2bJ
ca8sVYmJsUiWXOgbkoLGQY4KFxT6h2vABsIW41qBJ7DgAYS4hBhtkLfB7sxmtqSxl3SQ8Jdp9wZN
+uvOjOxl9L7Jd/LIsZ3PeV0H2Nu4OjizDPId5vtMuSQDySbQnmOdkTKow4StZbJtOPYRTdQFWcLm
EDqWGtYQeGKvxfFYa+7zYkH6jTxq1a4UwprIIjt8I4/G4SWpoV0dD/muRhA5BOjBK/GPQ+9OYtUv
Nv80Nd37uRudc25EkAfSGzR+vcFjfya0xuP1YsxVeG3aKtkYdnZuEgZZ6LKHVsQ2SqE6/Xf3YZUH
ar11WiT7LYPJVOO+8ZkH+KQN9qwuenCrKylHAaNqbAB+DUibyPTdcb17NHfUZTsNMDgNCLP0vl9f
Ze2t7wxTgEciwK99/O2zlsGov9rD2DhXGy1d/jyPpHVScMW1I6EmDRs4VMXG2jmttHA4xiYW6PX7
vdKTJ4nw17UW8ZaSliJ5C5tRY1v28olBTlO7WYh3tkGKqHx+3LspjFcMacp98EfOuWhzwhN5VcAt
tDoNHqNe+cRsPiDQC3Vcinm8N3Abg5XiqcTtRv7oxzNbk2NItKalhBSNgp9EjWpDLmq/vrGrB26q
sv6m8pr0VxvJVTsiZY98hnC6cUfQmtHtA7tEq4ZC1r81ZM1RGigYCmPhRyGcbJg9YGMXZYv0YT6S
l8l/5LlfsWMq7YHTMgipUVIzLADi4ttbKGA1U3KUlDMVE4Hiv5imKtHiysFo0vLDFTyRRDxIkfOy
iGmmZedeQ/o50J0ix8OZmx4GpZxZkFML/hYEx8FTNpP1U55rS0wYw53cMffUPUODHRe+ZLYk7HvE
0ZeYNQg5Z0Kn6K7nYRDBeeo7iKslgJqXbvtwe2VLMOVchT6bTvE84dxW2zxZXNY1q3qRMO84pixs
q60p5LuUsZFl+v3pGES6DCcYBYyr2WGgeoBuumCd+mHa8Prqdf2iFSXIOcbbLIWrwzAdxyomYTM6
dx+PVU4Hx0d2vPd18spddnR2irtLwxQq5gaUxfTY8pBpW6DhuwxvFw2DhgiH1/r+e4n5GqqRhydx
53DOM7fKTMpKQpAlVMmVh7dg9Z6Z2UowPr1LtyVJuqUrqkq5KMdaKbtZyQKStaL+nKpeupzUT5uA
EQRzguGACkzyjl3jANzdfOMikSXZ8Lz8Tk8oq/W7yvwhF2D7hLHRPLX1mvOOLrPv48/BDcOIID5A
ooaO5oDGm6QErOXD/aPil504j9afIuCVuqyyo5TKcBFg1M+vaP7a1QkZWhcMvbkcOcMxE2r7ACcM
vBZAkx7xScJDh4KErAqD/vinrBkcenW/nQXqEFT4PnAHq/7mzY0i73V2mzCcTH1mgt6KfAmEpe+V
3lpzHtiRpws4cwuprXanADF6s99/c1CV7HLVASJtlmp2yMN7Rt+Hefh8nzpPQFjNyUXKWdqduofF
hL8hqeEFSGXm4YIcVE8qIua4TpnGrvsnavzVXMZ4nT1HX5WNxaFbyGqmdzy/StY9SGZchg02a+UE
t8AaeuUQ8bhDuR3bjuzDIkWxb5yNlQtj34pZZ5e1QO67KPU0OUjakEuJ+p9ykfaHYsvKnVP9Vear
KUeQQ/j05KO4GhoRIZQsgpdWT1Ol2YcztgxRCfGSy++gUGSBNhoEM/DAtbqPX67XfpBP9hdV7jp0
gkp/VZgtDxgqXx0RIa4MwNq9PC10MyszBQaVY7G7UtVYi7V3w9Q9OmYeThecY/1WctEtaKZ1i0Kz
Hxmbo6xmU99A9YkAzBb+S8waqc+MgvRqnOJ7yNgd9723n667upiCucVpXXKpUf4LPbiezHXUHyes
XazK7TOgW+bV+24O3BZji5zf7qhdeFEtT4YpEIykTjlCmAVgB6YyPacdkl7fIoBY6EptXJc1DwJz
cBajJgVCQ35LCEGUkFXkNzg1HDb+cSraID7zDq3tnvoUylxfLog/IqCSr2Ksv2CEyT/P90+wkFXf
b3PkW/xD5srisraHT/bvUf79aV5tcuxjOI8G1+JPKAG5CUUwB+nyDlGMwpWTJHdBe+jJENRprCc0
usW/qxnc6JaIAZQlOwrMM16FRKR8iutk2u0vygpaZoq2Opw3dvVL0emyqZ7BluariobdPI+Z2kkP
/Sm1dA/2G2FaFhlSvr512ocr1KHf/fkMi/8CC4GOY4+VcTlRi+hcwK7QcPRvjNCh5s4xL0CcziNU
UbuGj+by2PzkgzCGKYLCAJZmLR3gH6D2BKgxZOUEpK2iY4QnJQbLsHbXAZOZ9HUm897d5b2cPDq/
e1boftCjLVKZhcfh1M5rLArebjfaIXJzY5xKToq96teITNSIZeko8uGl8MBZdcsz4f1ubCCnCO1T
2HgAZIxPSH4YC3K2PFVDGNOe2lPBq7vH39RDkIvj47GWQVduJ36fYrMvJa/DIvTccvmzj5/EPaYo
PVWCwmzg1L49SZgjU3K/bjzqyNbhENZ6B/t+Q3L8xIlHzxVLjdXqn8jhPFp4W2/rTZPBVmZAOSso
m+FFfRGr7B6JutAswDZFg0rsL3d42zj8+hAAfJpuRoYwjtKVDLWYPWex4rP4F64eNanKHw/IwgVS
7kRmmDKWcqJe0k51PqUWF0XexyEJyPCzhPZRfV+EGE5HRvmf/OQBlDqEPneDNRky66gLNGqGDRDv
zWsKIbS3NlG1JhHLsPNvdFpRkR5NWpVIujgI5Z9XWY2JDOUSZCnV93+4/F7N5bpAnmDpJjkS9sRN
sPcfsRQmVsOXT3J/+lKIISLHsD5YED/fUKf0RLvDP3POGEeAkiWnwbZM7TpUhPm+9LwvOpMBrGu4
M+5VFJCnHTRNh8t+ssdG9NlMmPBbsGXAixevaAoWNofkiTYBbSkkX023pmNLVKzQyWaxhqr/6x61
lNZ2q0R7UyEx2r1K7FKXGNRueNpxTz1l7iQ6i8ETTNVQjaZzME4SnW9zxvMWFNfOV9jzujGT2uZt
eZBoBwz/p+hCNhDa9BfjnR0VajQDRsbxpT+WNVEt/MnApLiaDYLLI4AML3m8Qk4vjE6jwYXoosZF
fpNt7ZFop2WvSQqYC0U+MJkjUaSmLdQFtGrELpzPaMxD+RjEPJRIIU1HxzERj7Lf/3Qorra+EsVI
cujL6tbPA1LBH1814usskvQr7cZbd2FEW5yc4YluH4IDs07TAeSTWWuFYc96Xzaa5BXemrUNQWzS
3yLE4HwExkXSVHAS1By5am6lX0w/fe4yy87GlwcGBwY+b32fm5n8YbXQgB2YRaH9qtYInzAt5uuw
/dee48jVx0sz87HzXUAfyEJMSTY/Uyc8dXnSX/ebuD9Zv0JAHlYYZh8bmxvUvzMjJiqVORZA/yE1
ZxLh1G5iyrXLtWropeStUTyTJhXoEHQtRumhj3xhFWXxc2kL09xWsswlGFMxX8jDYFB+GiT5NrmF
DgLNNADXxZZeW3tSqfKdMgcV+4wcp9kT5tvMLjV89oLfXDHu/4tuYSCsSKbObEsGLKKfScu3+eCw
kA38A9H5hybQsiXBzS1y1UXzmPYGhti1RhIzkwJwX4gX/Ar56Vz6pfYdN6SIT5NEMIY3kw4i2vC6
2z0FN3hAns3cgTCA4pU8srSzAZz4IMfSN2AQ4aKE5PURZ9ZdJjszQaZi20I2vaWDm/XB1oQ2rn6q
ihKyrilnJUztvZZuV0E62/zWShMpXA9wrA2FqBIDeyNZsQi2UKucUj+p6dZ0KMj+JLmaevZ4B+3R
ffGFa+3zsm/I1wLsUQvJjFn7pS+j172q4vk+p6jCME+ZsTykFlSKUHqCnAiJph0NmKnE0HY4jdQS
TzUrMIiLh6kp0YYJknP8crcERgz9MR2mI1swkwgrNaEYeh05qH35dG8A4oG9DbsYvNQ0abljOPOT
EysBHDW4xWSdvId2i9mdK8FO8aITKzMnHaIH9NnJz8QYIAxCuuDOXzQuahv50fRMKrEjhgZhHTr/
QX3n3xrtN3RDTSL5H9N4YOP6yMLsZaY32QALvXNXzikq7ywv6bQs0Ty6HYKq5ln4SxHXgpvgFy8w
31ycBUaPM3JwlbvyVXWlob1QFUWhZPuGa8Wt5UOMpfj3HBfeDlAFgp4jdXmnbdTv40gh6IHFiF2f
A5m72YZKLxV+E1/ci+39DpB0qUZRofwSY6lt0Su8haaTcIsG39fgsYo7y70H+YARNFCWtDq76rR/
LUt6GfoW3cmBmIpZqrCLonpoQczsm7oHsSVQiavxRKNrRiC16VtoW6ndLIuR9lniJjc8LsBz7m2n
F4m+/h2LeR6LnlyL6kuFpIxGww252jhllXQTbdeYODDukaosyl/FQV7AA+9xWcyQZ3Yhy/VnnChX
832CV5Eo5uds/4A/k6U+9aNdPWkpu0kyv3lhpqzYdx6PkO8yabtDdFAc/H1sPQz0ZB/6I02uW3+W
P7/v6iK9XQ8OJ2lutMSenA0cFlWohzkply6LusG0KG4178UjvUXygxf/JTS9fNx8A0AJrtvpZrPf
sOlM11e4SZeFRLBbRG5JMvrRX877h2TUc5c6hLmYmzXXv52Xrcu9Po4jdH1x82gYlR3p1P8QzrSs
mL5ZeSMpTnRBKIaRlbUWcUTa6IFpeYKzNlPKtjSJaOtKFZz1Esaafyag35uS88Nh8LltK7hdZ8KP
k+qR1L2KJ55ayMDNJzTVTHqVpmlm1XnlAeYDDkJ0uTjkx6g/0ekZdx8hfABlQz1pU9toYTJa7Wk2
McHysvNOO8ND0BJTZJtmEfkndJ1JirWoBjRspVCXhbjC+Uul1qAFUrzk6nUGSqZ9JDWqPnwHp3I5
VuQOpNSachs0/fl+TipR3U4qywC6iCKGfkl4K0iPg/o4/KAt+fluffQnfAvPw65r9VMc6pwVh2SL
jkbIUH5ZpWdHM+qa8gAL17diRaaSF1WDY+gK0/pB1bMIrJ/H5eozElDm79hHaWyxc+nW22B9vtt8
YgVoJ4S+n3NOZR5z2bQSUUu9YdDCMaHBkq8yb0wcrXugiGb/tFPzc9qBVj2xZ57avkGnpmLgyQ8r
RqdDcfhrdsmfmR1nP3tRcGPma+OchrfDcxtBUTBx59XHQ95QqlJwtrCkbIDTrDa3+T7Jh95UPw6U
mZgWUXzEFZec0qyNchgXerPiqvKTI+7wnvKeJplXe9NeUqFqHRPf2TbsyTp1Sz3H45SUcdXYSxh4
2FlOeChj3kYL062cnUg6Y9lJ4ooAPX3MBAoE78CrQPrGfq/KziiyjieMlnt46Iz0Plk2mObqdnix
j3RBWGX/K6fnc0K9KDXScRLPfHZUpQBZVjzNogsaKD2giaZ5Qa+O5lgZ7mzSzPrNyAvwBfk4/Ujp
gAT4n0KNyTm7aVNJ9JKmNF7mVd2wWbLnF8w7NiEAAeQ3F/GMMfieN97QjAXSmCIpN0S5fU3kDjls
Efrc1ebxNU01Fe+wTE3RNIRn7RJezXuk/mgxZ/Uo7/5Dit3VaIrK5q/rEg4SVRlHLRGrS9op7r45
Wh2WZhKntmeKXn4UeM/qFXN2RbrJQ1oA5U04sPRZFo/k2g0i+2392cKmpF1trpZ9PQ/9aOjh9OiY
EkHFXLscmm+yicABaxzuhu+4Fp4kwABhJp4mTl0pt4d1lJgxMLlTnGFUS5aD3BU9CrE5yk5pKNLN
duDR3LYpgh7pSyDc5lNv51pXL689oeSiqV5TBshvghoMx4s8jSmYIA5nt+qA25RCM8nWocC9jc/f
dKXi0cnQrY8k0R8WP7Iu6pUztBqmKFf34+epb2EBnoWA1spB22GE1T54p+DMkyGtCRtLyX5U52sF
jArKBC8V5ZnBljoX0erAhXGImX+hGX0TAmcVFioxljrPQfP0hmjGcLmrijbzjj6+ePrXinsfjKDP
tuwU5qmeFxPeVOOMqaO51ECjdhWkZUV8tDUxLJeoEoSSCYYgEL/orX6rd3WYLyWPUv7RBxKd2alD
aX4IsdKO7wlX4qFfhsFdTAKEXnsSIH/v7dYCiZOZTyiSfbvD+rsqD+HBb4EVlETb9m98HqYB9OKp
AuwJ6rxpBCzCCnRj6ZJM4Yzzmjy7K5JlcKJVR05VFTC6aZu+ojxsFDgGzfp5DXhO+N5Ha9QsY+LN
wGHY4jA1KmG6y07LZ8PrhXqfIrnSk6V0fKQ+QlTyYd4jaQ+zSjpTV3VPQLJmJuayXybV6bIJt/zE
yvBhF76snUsNd97Wcdz/ttEmWqYWiXJGWEvx9/qnLSK9bsmivDFpjC8A/2X1itZ/rhxtHvtpqC2N
NNVBdjFEbXbEltUHBnsGsgr0vPrC9niSIRFrUS5QCICZYFSTEr/fS5neDC/nCSwIC+VWDo3XxRtj
QPLsN1D1OFA53zCyd2hMzU+twKXNYLfajNG2WKbKPGqHSocg/G7wUR8VAhNbYuQdw+2mQR80czxM
+2rVzvyus9W/RGXsNCD7+mdTfTe+2TlgQTsB8uRZO0A4wM4hS1cfEazIKtMxB2Odbpt0oi+JMO4T
rezIUCEL61/SNty8UtRpSjtXulNUyb4pgodUb/TFk/hVTiGfGx1OUnpkwiHuSogA8u1CHkOi92RU
Llk4OmHQySHzHKnuUyy9owNLzh7iATjBNqm+bG3FPL6iY2qjyr1d7laVN/09bXdRz4cuz9BJdE71
n4JlWA9SnE1OT6E8nJglRKEL46t0819qxLhcIjUi+blpFUueqMbiSIhcdDh2iuyEq272KeMmmm77
jwdEqyS4IrEozGABeB4h/FKw3/iYG/wNxRTIWtko6unvrCPqYumpgY+S/BlagCQrS7Ayy9uXIQjy
n5g6rAjafjXEAev/rn2larws0EfuOyr1IZuZgn6N5hakE+HRq68Gqjai3XO+WhZgZQk+gPhBgWdK
ctr8/AKQyvvLZp3ay9xcdh6I/9AybqFopWYjOk9QpgGaE+2VFOsgrZSvr1+VFS1E0RnyiZrk+Izo
P/pcd8SZOcKYJGp+YcKbzYSednzuE1ZX583/JyxH57y6ZL8auY7azs4JRhsFMyB57FviTDXoL8DM
zxbsdPnICfiqD28T1z4hpSPrTyq+ItiWOKs/7NQO9eOikvIEg1XN3AG4us5QOn0OIwKo1NtFrOME
6nY7Zj7KTc8z/Ovw46SibfL0cLCQssggnMiccOgnTBU061PARQyDW/RQxw193lvthRYm1uMponiI
JSOev+vU8W9bKhgiqRhZA4PoUBCophXUXInZ3cREQi8kMmLZqmJmfZHDjdNntMdtNy3zDLKoREID
fxoDchB8RZzvyCctqAcItoDe9BRi5w4KncR8lCUh3Gi13PSng25N8NNC83YBlQxkZQoXlSnsac2f
BUu7EMsuUAE06bn1agOaYyAc5cSQx6U3cj54nqwTHYrFpnu8K7u+KJxH8WZkkX56bmiPMOwtbxDQ
LoKHhoQqwl8Y0z0ykoakh0Mm3xqAfV+7U0o0DdNbNEMXztAN+slrZ9ZnLVVnKcQjfoUOAo6tzoRJ
+olao4HjhqdxWQpIVkE0tlcYlW2XwSx9EUddgI8ApB6aLg2qudCEHZHv1EiEMBc9vAypHfVDJizR
Iu2qA1ZIEdys/kU4WSk9MUohrkXS6rmWjpDdwOlqO1n4Ew8rCZ1jEDWSuLb/9Mrwa+MDNG3tNVJH
hM9NytnO/s4ywzfk/RFa17RThS+OeBFE2GzDoLOR+6DH51rKdmk/pvoTWr0/G9BUrB7F4+EgSoy1
avYLmxCAYBgdFGwNqmCpPk5wqIu1dWnic5pe6UmX186H4ZKejEvtfGn5bobFMB1/CatKMKXDigHR
aNIafZAjt7E3rMKU5UkmtQofv9Y/6y7QQg7kat2PCAZPZLYfa4brg4poJOC2RHfHwmRZokCdyEAd
dqKMnFIamaeTUo1L2h2THxVJyZhjjkG0V7/T4Cat2t03+ouU2JbLz3O7kUCTDGKGwIzyI/nTYIuM
rHnvynWYw/3ETdpP0HZPNfWwseEIGq732mP2+H7VxnO2AASIxljGDXwJ03G0sveV0oFPSrQ6bWaS
mdb48KtipNibHZvxwYBt5DQ1dv4nF2dKz+YBwZDaed/adtnVTgIzGpwuhiR7p3jaInG4hPJeH28f
mQUvwT3NdLiYP3Q8Mcds6LTQ1zcZpM21RwrpYYDvA7qmP+QSoZIMcyeffHSCCVWetshKNH5kBCvR
VqvJaExqJBJf60xMvbG9q+1ZHfn5iWqSrAYUqY+YINpI3XqvIMT/Qlz8K97zl2EmcFzHqSJbHKur
aYJh3M0FKf0sRbBartgUV0eiHO5NfAebaplS3l0VEOkaqrIQqt1jV740oHkGl0xy98hcR8A8UFH0
jArbWcGc9erotnbrqt4aMCFPlSjdZkrCO0TldKT3O74JlwKPr/NwWzSDRQS4x8YA2PYMC6I/ziOV
0XMADPWHMNWePeC3JMrFdonc/MjzGDCqVZ2dOmaWr2Wxa8qJTylTNYrdBQS82uF9KEyGh3vHZtgQ
AA481XrQvJdGgdsaKgtsjKnDwBTTuV7g8xdIUwsERxWnBuZar0iYialY13evNM8C3gql82r/fJgr
ulNaWXpLAskcnqwzAKhvYE/MFGjPXDZs2EqhNSOkbefJq+3f5olh16FyzTJ6OwQaVKxqOAne2+pn
cbYWOvQM2HRZfhtlVzDxx7cg7wyjgOCuA1uU4S1jlXsVpoaMu7SVeoOYRpr7nM6Sf+hGNKixOA1r
3q82OEQLEg3549Dsf4KM0ZFrrU8R4HLTv7VlBuMOT6gPimTwk9L0YAn+S30S+BUMZmvWQNalrD3I
Bt0wyhY/Pk3jxLVjHHfNDotLs0H8FV+fdoCgvQJvB4SK2tukHaa07mGpDMEl6avvGp/iE6TBwWwX
kF34SB3jHNMtrdGtvyQKpmX54Gbg0yiVRy7pLt+zXHEIdeiEToLMa8OB57RI8YuauQL9zi5m860D
g5HXB/wxAwDEPai2KhqdNwCkLzl5VSzCHKrNL6nCti5q8aQ+Ru5LNtS4N31ChfPCupIpEP7ExM2F
Qpp2PrmMUknZI0mXCiDYh9xP9gnTMKqUxzgYghZpCgCXIEl9/gik87DCVDZkrSCrlaG+ohurKM0+
oxWN2u806jRexXyikDtnmfOUgHhQgDc5Ox8Z+M3xsCxpmre/iKTkkUvRV5hRVBiCLOdCvFLyAOEo
xuzMx/WhroiVpDQwPR20DNSqNvunojhMBf+0fJPY+/2AXcQwtW54cocsHEpl2r6pWJJa0mtDbcyJ
Air+kE0jPLSbmWCsr0WiXd+Pp0HMwEol6hKxx3mrjYT0s32kblH0mT01D42fS9vsrS00WpiAOUTB
vLkukkX6NUhrcIqdQzIYrYtdLRDIj8hxLaGukswYPgyKP6s99D3dbXnAlh7eR25AfiiuqCbdWXJn
rGUCrHmCaogasB0SN2Ji9vnY/MqQibfptBRg/05IHs7ohMIKlawfavNI+0yo8ziOrSKBfov/SCAF
Fl310GWFXdSWcs0j8Lx+ig9KONZy6mmIFjl0hF1kDsb+wuoffFc3rK6s+Ufn8kSge5tFd7DCYjii
0558eu3OgV8xc3ZO9xdw/yCoVRnuNcRvqXFZ4xWBFgdRz3FKRqfgKZUUlfH92LdZaqvdGymW3uhs
zQoTCF/F6RPzJQu/+YQVJMj3JFMhfa8BGeK4ytWD9TGnYk+FcqkT8e90i9hkwU6s56IueXxJC288
yLvWh//+F0RBvBfNyk94s8SwF3qJ2qoiXT/5rB/ZSrsCHhz8JmXW/ZAsRjtr9t/aSm1s0unEz2Bq
YJUVOfv5el1VGo/rMWjpMVIE2IMxAuvidegLabeDubUppbjuiCM/DBZq8ZmF7ile3YwoFw4cmgiK
5RClTBSGzW/V4Dr2ACvzzt4BxZ616DEnyEnuLkum03s/cz4JFwBXa8mFQrsgVp/vqMYzBflSWGlz
W4lMDT/vSOiumLkYoVoXSym2jbjAn3jaZa0YKIkma32dxQk8tvD54Mj3BTBiCxF9nqEBqwfqInXP
mw52qGnU7B6VcgmajBHA6J4yrIkjzlvdV0jNrfNsppMeJCaKQT/JdNPAqLys4S7IaIOvaVFLiWaX
+Bx67cA7SjUK2OkOrAn2/8jIx+EaW1xiIEuuvfg9QVUs18oDRZzDPWZYNaADeo4wgbxII/zEPEOJ
Dc4Sbs8mfSx2PetkVSw6fFIXMUaV42fwMnevx0IJ3k4vU40PpNUNd6t243LhjgclvgznmziCPbKb
CGZU1o+XHTYrqxgaOn/qmCf6gYCPmy0Ws50G0cfF9DDD3yMQtzXJP8iCXFe2mDpYcQFMPqNKYTlG
4Dr01bgtG7ek00Gk/S57eCQFSvH9ZybpUcVg+iWNlo4IzRhPZgA0M0ZEcQBitrEclMZNM1pLfrH7
wp6Z0u+3V6k5bBmCkOIDDkPlTvKpTRNPW0IcQX7IBbgutOBp5WO4PKJodpC+DI5NNyzF0sXXbkvP
FfxW9yDGwyStjf6dKd2wMq1sYDcNCi9nh2gso1gChDGJUnGMCsVRCDLwkr6sKQdxLXgR5K+fqCDA
/BpzikVEZGfgJqnj97EAJE0G2EGhhzqsDTDxvYtH28H3Ti6KIp3vXTnw3ARjXjyF9DpOhmAul251
N7MgccqWXWaeSyVo6nsrHxH9doxRm94ru/zqKSlWkbsG2l0fnp+2twj7ssmB0fczYfdPqwcfI/wh
tl0x5nGLXcKJvIfyiZOw2RQPvZ30p2x4wBHqm3yTPzFPf0qgbRudRCjV+c+RMGN/yrk18ZQa8OQb
t34Pxs9xnrYYS5GRvwhJ6AlpEXCYsCoJlnd+HzmyJUNnrM8cKxSEmXJ2Bq3YnNkSotKOKrazvEsV
hqhXTSCsOMTv/HauB20HlOpo5ZA3QaH0hkx0vA3IHXVnIzbSBQNxLoxnm1YWpQbbUBouDxXlcaA8
koXhIxx4LQxH3BqNwp/DvqHpwPnxbwB3fpACORWxLEP3ZKS30BNbXc11Y/k9C4BjA6VCc7lySChR
fxa001wfTMSWoAR0SyM7qhpDJQRWb2W4bXA6PiEm3r3eJ55GLEhVXbSJ16nApDv6Ce59i+5Noi9O
2A258fTBI7Gi+iSwJBxtS28sdtmPwOHq//DhjiQKyMD+Hq6h/WozGNkdhR4YXm/o/j6rF5fAPP+0
vv2iqx/TpOKocksp+hz0+b/ajTF09TwEthJ2Mb5w6tHKqc/urAnwkqbD9sp5yQFEAg/5EZeXBnks
ca5ys0MtNlOQv2QPiOgEkgFZHragd6wwjE7TtC+DAnqnYoW64M/GgF39TO3fsczb5TOkbQYHtuD+
lxdXd6NpZmWQfpVbyZjv2O9wtZ+LrSc4C6M1jRQ0Pq3+XarGfBcLZRBCCOBmvE+rQL79cZ96VpdF
xEN1pNRJuVcuGvpvluifZEfJ+JC4YYYo2yLeSCaEiEIIrod64CBDb1XqkS0RC5BlleB4ccXjfsZO
lJNHe4qUjvyrjz6BrJv9I/2mghcjj8QTA/JoNKDnGK4fQc4VULYhTST6vRf+6d+YpuY8sSgYKsoe
QTxNW3MGb5KYfIgK+OJHkWQXHHG98jCBls6EICcLiSFAeSu7/IRDGrtdOYz7qbWkhXpU29OUxQvL
+CMa4nbvRwbEZgIwGESGZ3UQNn5rb3hrtrSx4UYCjA1eXwjc3ZF+uEVe6Y8d/+3NvJo583fXqzlM
L+osOChTsrMTufK9nY+1D3SQxYYiwsknaTY1iEuUjhHwOrXi8lUtz/ELb2lI027Dv0hHY9k0UUVv
1HwIUilX14T33IIvMyWlz3KBVqnJ4dodw/dAaNqXgNFXV54htj6rgw1FIeAG1sbGqZhgTSlyRaM2
4MuBZdFwStwQIqk/iNt3K/UAVYuMOveHh3E3iyUgo2+Djb+5eDQ/XBsbo39zp2iK8Iprn00sOu+Q
WLfcgLO7ZA/7HIv8Pk+XOuzR3AsqvyAGBmjW2jNkSvKAtnrmp4pmsFNpkMyJ88AEr3ik7eaTc05f
pXg/S13LV9SeeIw/cXDp2rUVlCUnpdE/w1U3Iz+Nf6L8n6CVUUtqsnuO6bWzqNz6rmTgcWa+ohp/
sla2vPb1gyt940h+64ff9dvjRVaX7nkwSWj1frpvmHTvwvas5tmNelLo/4JQ5GOveAH2Hl6A8+uk
w8hTso/HkVgSoGkQp9h5W+baQQ22OliroWah8lNg23VD9oH9Xrjp2TGAFxw8Ddju1L8/P827qIve
JDhtqR0cZBeKrBzzBbN20maGlBhilDhWz9/GNwZpMj5PjDiq26+r8u2zFyJCH5uYF1B+2mFpj82A
ruk67wq+vcGRMYTE7nTLIiS9vcnQzc05lT+cN3sjKJVIwLeMC3N1o1sAmk5HKAP+4K9MywISQEJZ
DFZbU77z9gevsSvXWPrFqztpV2YJOTef26zWmdSBhlVoLheqD+ERcVTPYxOCQF7ZAqvsf0nWOkPL
EOIW/3j5H0wrawpVBfOU44+5u9HiCw6qXCKiKuxzHHL54VSnsY2zNUYw5pD5vNoxYX1n3AmcABcA
5RdPdPUzgA4JJ55JzhPQZAVSsMrG5Sylk19RE6DDaqJLDkjYidB+JmK8nOApsUoVdBqb6KU6BIR5
l5AboZ5wCKPU2AVdLI5nyr7v+zE0h1Y6cA04z8YzEBBr6ydfSd2982TeAfRQuKqENGss3mtWeDaa
RVdbIITpTieNCQFaWS6r3X0TAK6NKHAJ31SzgaQKSew/1X7AcewwHmqw9TEPihs1XOV8owuOpWB+
gtJgsq8/E4Q0vGocZQqHmbpMVxMPGUtHZjMAbP2f31Fjj+3uQPwZt7G0AfZ60egR4gGX8Pd5miDC
l2dYHw5IRJ58fVdHMAe1UUObqghkBhMGC1Vs2/Yv2T3F8NnYAJ1HZ+HK6OozNXaiS58dbbO54xrA
UPEaUdmHPoWfZ2DCDBbDJu96p65JYuvjT7hcX85xx+Pr6vm0Zlg/fjOQPqN5GYpRF09wJgBVzH9N
v73XIyEPzYAPgWwu0vl9C4us/TvGJtPf+OEL5F+uMNF9jrqBiZbJaulugNeN8MXAM16J2nzFzehH
wlapJ5630a+1Qki6Q91f6Cp8mWYRqS9kEo9qq2uJtWjF3i1+TS8GMfcZwdeQbMHxk1u8BpP7G99d
x5BSdy5BfzX2cDkPaEnDs3+Y5kHlSRs1eWB1SB41QLFaV3mvieZfGKcBlqjKJ4FLVwwZ7zTCnz1q
eGO4pwCERAIB1H3B4LdMBbViKsEe8LPCGjF21YdjtaitgxZgDLPRuOIHb8EWofFXrykLpeI9xXuc
KW71GdRM57DAs1krqxS6CWLCtKDJJD8nmORrUUdknzA3MDOjU7S8gM3JENUa4K+6etMSy8EbykU8
TyqcDODoshljPJipMHzRA4RGd0XfgVmbhaRSH9rFTVlX255dT+J0ZROG5lpUgZo89JryZrf5EJ8j
z7vImFfFV65cqjttJbXBTh32a8tbH1ocf7bh7eMWrCYclKue8thvIovak8KXe2RZB+PmkUzH4DpL
OX3Llx0/aqZoObxkEA6uSqj4WjWbTkK9/vBkzH3uXBBRIZiQCiZRlvbEcCQPasx2ySNm/zkuLZs4
Xln4Z0tzK8N3w9fTh790ogF5e/S4qRN8UiwpaajFSGUiIeXRx3gf2CXl+FP6hHHtoytB0fut5t/k
Ba/89pkbFSLIBg8hM/1ykvcnZSEaSiui6Oaaiydpy088ALAw/1xR1X0i1P2mUDwmpeS7+nRc/P60
zdzW7kL8tQGKR9zF1inxgnIC2wT+FEBx3bCHpF1rm2BOytLrRrI9ADB2uP148O7VgxZSVCy46iY7
3L9zDXsbPC0T5ORKlkhx9/gKaDa3vQPFz0Wugv6QxHerkdRI6lnXJoIzJm8Nxwr/LwVATtv7IUkL
QbsZuNMSrmESsKpVzKje0m+4SCYJioBH9SKPbMfrTBQFVaw3uu2ntcjP/Ti5yHH5kiG/kHaoxAZi
Q+Xiq2uu88zto4SyqyJUDn9Fanb9PPr7b7FgmhMT5dL912auTYqNmSgn1eIuAsWkFMxH5Y9pffEV
xw+6TV0oy4SwWsJWI220J7A0TK5PflC0mtB/j4DYzbduCFNXcqYcl9XqtJxEMzRhZxBHLrBHWAY+
ObcbO1ZNmdvz26LJlQ6RpmgEbOnuUaViMcvpV9YKN/aB9LP8k7dj4ZEF/KEeByRkB6xZtWLWhfpD
Qri9wjl15C7OWR+UXsN7JUXjrdhiHVmVQBh62o8XZILSzq9qkLB6hAS+9XXPlLjuDPUJyWAo/DYM
asWfT0OTZpZHveFGiNrzim8MODZAyjm9A8DsiUx9k3ugn7KyQkpsoINnZ+mL7DfdW0mfIJBYC9az
RSlEzoZkeNGaI2N/3BuwnLDU7JGnUTXp7hzyuiwmn7sAn1byGpCKgZicDzQaktuxK8ywg+TfGL2T
PShwgD4/sxUQX2An7NtoNynMDhHUtvxvLPadwd8Y1Dp8zGXI2VqXkKbqJkK99bY1sqg3a+Kz7MSb
p5jYs+3ISSNZPsYz7aGtPw4qPDVKzIbPIm9pUagnv65mPNoTI57kirHV/zEKDCxOZtQJz1BGRNuq
ibSKcbSmx6w/qtRm9PasEVTzON3IxiKhfzZwnq+k14T09uzaoJA/RbVyYX6jXPKqyRzZyy0EdO5n
t2lwwSI4JCTq60gNXxcAZ+C3vCcNW8bx4SIjYzPqTVZ6FilJmDBwPSCL62CFJAk2Y+G6NpWf8K1+
ZCn6KFXCltUnEB89OdCbukrZX6EOOyoBMmXNZ3q8xzkGdz7vcKzQRbDwSS9MTRE08RtL6LmABcIY
vTqBYgRbOvrWt8QgdQ96hYJNdSUiosBvA+MC0xebAQ6BgfI9tZghlibtw42o3KnDWhRDl5jh+Alc
vtWC2cFSr6KN9EIPEns28UFNLvHVK+3aWaj0r/ftuG1wSh3xZl15tmD5L7gM8fttxskz0fcoA8ni
N1pExWaCXpRVtHZOohdVZv8ro8cty03gW7qNObyJBduktPSD7/EsXV5LF12Mu0c91e+Dv9Uy7E1F
BuyUwiiR+zVwFDZ/M6mBZpZzhFQht+QT+h2TLR19WdXynB/v/U2YX5X9m6NnA0P6KyyM8q5NwRi/
D5KCTPKorprd26LSL7MgrRt2NXg/bc/F3n72yWcm39VRI0wdUCJgxSRNZRj82upAEK6jeOFmok+Y
XKZVuqR3tI7uqh4+4aY+5LErW4/ixjGjXcNatMVbh9JXfXHHZHnGpQpB4XR7x1Y+IIJI8NwSt9kw
kmD/6Yyprto5HT4vG5Og7XFg/pU9vbRfvxiGy2enHl14ttxS7jNpWnocBlEWc35HGVTewKPHhAo9
Ozk5FnCX4SD1dr8aEOp3qGVSKfcUmzLcqoHuvkjA3JPTyTaAemCw6Iyz3nhx/Uj0e6O8Ljbov6fD
qD32lM8BjGMcv7rEfZUmDWL6jLV8swZ6mhsqJ5Dc7GyjviSTxXMkcEFdgjlMH4LLWW6GrKYsugb+
4Bnvd8iYS0zHqv8PSZB/kZjjtH1VPy44UzUq6A1X+bIZMkJHirP+dy55qYsKlQ0RI6VhhARri2v3
EWqjvlVPGEQFiipCuw+L1/j/oUUgP0ELHBaZoSeJ234Ju09N8NhqS8DVN/U8YTicCGapNMViWm5w
LMxJh5XW4WhXJGdRpIf58SHNbOy88ftnmJTszfMwgVbxwo/N5xu1SdZo7L0hFk/F7Wvklaibj7bW
M1qv3JxRxgN6HqGZj5gsyhvFyNHF1ufgnsSiXryg2YSMq2TxOtsTij9Vp4Lz3+rmFxMFtNUHyNb7
sFixjgVpClPGU4nV2B/3ffLQxaXjPZ/R0FvFFOdqmsZ1ITxI0/ox1hqFJMHEI0j+703qov/pOlPx
MgLppIVJgqfpP2Rq8Q8fvxvdvgCyd8bz3RdE060RVbOB4IcUOtJqsMCZ1LweC0dfCRJa+7DrkvO2
IBexH/QBkmD3oQ2h5V1eIN4PVCoDNQXdRi5KjCtrfQT6l6DNNnTrIOhDnBu3RB74eEHd9Qc2/dty
odNXEqpBvI2Bz19sfDR7PF0Aa1XpMorBM0nP3pNdcK3DaifqcNMzyheb/JAS0z9zZFwI10XnSt7C
52dM0oX4E5aiIfdIKDQxSNXJfIDUU+X2AzXsEhwVYqEwx4VThSCzQV1fH0ROTMxrfw5fVvZooxXc
s1qhj1fhneLi3QQO413LlrE4ajqRWNAQ8v4HB0x+QjqPjgccK8l3FZdnmMeUNLO+2SgCITWCfb7F
4akY84NyjWb/KZDdSs9lezNmHKvMxagc2tNSz/5/AoLUDtK6aYqUiLNudZuVtcuG4NzmLszWjlX8
nyknWKYdVSM1YAjv3xlmvAw9LV+KSq8PRPr1/KATL6OC9WNgJxUnmUWMGDIHDClNItQLR2ir2Fg4
ABws5suZ+l4+5DIb35daBNX9zB277RVcFMofRdMMt5z68q5yyTps1UlkFJguVeFo3JLv1S7tlm0t
CH4oPHPGlzPZQLCGaw6LCm7hrMm2WaK7ObCFc4qQgca3AMfA+qPieHDJpJrdJ5iL6v4MSwJXvE9H
v4pOsL3KwV/VB883y2s8XIuuC/I0UEbEiVT6Fcrtk4beNdJGUgLUCswXaM9zIMXVGHV59wwNDzc9
80iABf+Kcjvz6hjFfjjIL53Dr/YNl9CJ4QaCQzR1XuAeZP4zP3UICeertkvOC0cCiAdaAw4rMw+9
KZDsVDSyHQBCgMDxb5GU5e68qFBFzfaPwRZ3VQFx1+D89rEC6OMekZ/GiqBG/vdBz1GH2V95oHgp
mEarhdiXpL4QB+1+r6TynpOF8EfEw2lM8t8s/LBtyFZiiMxDwwdlRP16PHzi6BQsn9iD+//0hzda
Vu8ua5tl+4uM5moyXWoRpL1rnlqCCuqccWOgPK5/2jzZoa7PX+bW4ut67DQ6jGF2m+0dDw8ZndPc
8cdaeTR4aQaC7tj5WEYxVo17+uQAn7KPQfezlYtCf7CF0gAANCCOGhHriR6U52kCxaM4xeGj7Mgt
114pmEDcukOdU4kx7Pka75R5MRBiu0WCAHkFLYBMV22ZG6tikd5DKGCmaeJ0/jvIMDpB0r6FFf5w
c/XaqsyVIUio6VqpKyKIgCA4zm0RrBxrhMT3LGM+xTAlqBEKwLOb/Mj7MfcXO1bLcyKkLM/kD6ug
bhm6dhTUr2DMM8wRA9H78mLs3ovFp1fg/MEEmY+gchOzvaKsKp9ENXubjcoo4tLzgwv5uz+ozt38
FmwzlGlL7LdOxAjq3G5NjLwe+zYhvUM2+VC6o+K7Kwq0JFVm9AD9V5CYn1vkfVeeLwazQwVuTC2w
zRA1n6Kr8cxpQ+xGjf33YLDhHg5jUZcxvdvd8zo2iep79PEHUHNaPGaJudzlP0kFpj5/8+gHPPkC
oWj3ACnRKmX6i5yHT2QzLyP0pitF3lhGHGEiAaUxVT12N3TZp92V+S8U+4VvTNy10C5siBNcVZOQ
/sonzfoaGQ1sctb72gNJrd3DACt67+vfaM1ckTeXXl7dX0Hgr0X0eVNFLONKh/zbrDYQ5+LL88ei
B9eiIONKE4LWFQTvVJ4D79N3QBNtdE8jPB7K209c6AHuy/D1n+ePfBXcRyGNvdsHm+Mi3ovTTRZp
VfXucJwzgY7EIyN3k2P5IuLKXtwl3qZ8NGK5zZlFyvPv9NmqPtCa1jtBBfsvClAfE1d6XtM+61Is
YDdXGt6Vcrv9hZS2+AK3/57SJmg0gwpR7WFDrCXYLFc0HOts5uwggQl4jQfcRAbGUqLnUl03nSzi
5X4cuxvIOmMymuY28dC5FM8yFFLLOsmsosHJH4nl0V2Uv0jEXiuPHu00ulJg1VWjXKbgmO1a+gPN
At+yHc33i0rOm9mN/CJmUZkhdqgMBfxYxKDNvna+oYPb6AArwyDyC+KpSK8In6UDA2w5yfCvs59+
Pb6+/hvFI2q2aqSUVAskM9FImYAKswaizr8xLD7zM3LtUhQWwjqPIPXcYqS85uSKhif/boSIt/y1
88MovO1HJwvloitskM3PVfhHxHePI/gjp+rFPXb96qDUk+JweVTt0efHlc65K6OhGG+eArYfLfnJ
NjK7FwCBVyvjj8Vrk/Cr6RxH/OoIzL6e0fVvr+DieqBeD4/fk7AzAtixXnGnsBlDTK+XMBE+Cnhb
0AzogeFvKFcDj9TKAzLm8QbL77C+r1p6X+mMHxMfAkh1LIEJ0qM5njqOE23yyrjCPO7aPV0rfo26
C2uE+H+cLCJKGEmblJA+3vV6Rbpah75sSqyd7ClR2aGoQ9Vksj6K1HdtIZ2xnHB2GvncwAt6yp0t
/vzJeDwTzQK2LUMGfrfAANVq1QCl3zvpJ/Lsk6OcVqN1yklnKK5iFaJLzyNybnltjYxAXpcxFhW1
pCrtPPLkHqHWwAyCOSbtR5n724zDzG8Xf70J/lgutHZVgyU5/56XUMJ8DMsoVspSgiVRBSSZOZ/7
6Z09DIfRECanikDVY5RYNCHRB62cOzwhQFasrH3ekTj2LgpbSAtGpBOg/3Q9IEMVWiAYbX8/RDhN
ZIFkdPjFBixAer44tWu/nKhnjbGC9hxuz25ap5RIFXR+Ij54SoFeRWolUPam995QnMQAzFFL9gHu
ZTNHXz4G5gcsJaT2sx/1ESAb01fHtk4xUc00cZFaasulUWZElYf+++7oIymSE/tqUdFML3edXpeJ
Mpj2FdX415+7HM5p5Sfc77IhUpA9AAtEQlDk5EWB90e24ZptybzvyB0onWZyoWv5NMdSTL+I4mp+
h/UGps39wWRG0CT8J0TjbxrbPw3GR8Zanba9n1zrLzvb6ORXQYSpWM7f7mZ6uDkGFMrtjKqS99Sl
PNig3ysmAtaJOEjoF5WQNQhwceuU8KBNdSppLImeslIcPe4P413DYf38UXKv7jx4poC24m9wVH1O
7HkMTC2sT2bIdCgdH6L//qfzLr0yS+P16yLEGT1UklFB7adWxJEAq1WlDCsql/9cjkYHIwV3Cf6k
GWXfsCinp7S9NMcZzlBT464OVrx7G5Y4m0/PlVrhMJtIoNSs4YRWsKcwxX4DAATcUmpoi7InsHR5
hRavaCJGegfq86s7A+z2bCJlzEfqGwYGrB/2cqFlM4+WK8Lx2CJZ+k9muLK0cr46w4r7+LOL5Uep
a436XkQ77WEbxr9tbh2Omh7QL5ATrp9Lx7y1EgMNKw3FmAWLEUUSWWuLWKmRVtellKP5J8Dalbwb
6keEoeB0BbxPmZ3Foqf14MNcUDZ6hNcjEQs2IzThPytAtr7lEPIQW2DvF61V5gTlg6E/adb7HPCP
j9N5gPg+qRcvxaqpVHVWluF5DlJkJyyeUv10o1VxJRedat8SFXOySnJg107WaFoS0fg64vD+aIU2
Pz5LFcH5Udm1hxfd9QuTozcg2iuygV2srGVtQeKxwLM6FaeJ8ctgh3llDtdb57qfOxksDEAYH+Y2
7JEcoWESBOaQEINxKYli4vYVeyp4xuFyU9cnOTjxV5oavInbP+el9zm7aEpxu97kSs6UNzdVYAHX
qYfj34rJ8QHzaG8qoS3zXZyCimKYyzDj6nqe8CtcfiiDsEaIelZhLQ7szPqK3NcpZ1+Q8nNVQCQM
cBf2wjkaFxdRgZk4kuR3eBBaXM5rN0Lvh8niS9IIkmyCrw/GZLhBJ/sm5KDaLgM1YejWneRTVHCd
7bStv6YUvsS5z3bb4MdkNn2JV1m316iRc8kNJarUbuRGrj4C5L7v+ds3kqxjE2y+H2jSR82r6jzy
vWOvD98VwPYB/NMQOCWg44D6eu5AFDfy162apc9fmZ5zKi7mmil9OL8y7KnHqFV7HcHmFElzIjAS
wPW/zhTClILmqszECAhFzrnqcMYmopvbutuD/oPLmgpYP7d5yJu+WMCI8MODDPWE2uftm8MQL3ch
jYjcAvfjfwvgXkEc4ifiqIP+ntnBb6MH/qIjwcxrfcG486/PirYuC0qSQ74Gdr+CUIZw1oCIeoG3
gNYcaMe/yrnRmwv5peJO3z1wjPEBcv+5HfYaX4Yc1JQRfn/WlwvwwspwQnxon6LHWKdP+9GAFk9V
RWi37TcLEu0n2RmJxSd4j6OvIHX00YNnda5ziWCYvw2ft68VGzgAVlw7wHFrLNlt3nE+eOFrWTiD
hroI8d9krOWHwi69gFkgWbVPzeknZpK+rI40KhaVR0+0fCugkA8xtK+DpEGclfHDMX+E4+GFRPtp
y1ShyIRQeLuxN5eKVWj+G/H4oH81A+blw8K01GfzML2sOfRrZwt/6skJ+eKFjLIeQ3yLpni5LOOe
bcJjpKXnETW2ruCX9fc34jG+SQtvyC/WB1ABuB+5FMPNj8gpJ+si/2bQ3B02ZkYlXUMlUudrym5d
Gblce6ee8Vja+8E7xJt62W/7ayfHGpKNsEf7W1RQrjFwiC7QpET83RtUM3FHOXVMydyDd0PklrYC
CJpKVcZdyapNIc8mqLf0eEPW4+5pW972RPhkuw3NSExAKqETwYu8zc57gF7nNye2ot6q+k5JLS81
kOkJIfNeSGxkKQpQE3mOuJkAXKA5oTVc75EoVtU9gMKonq6I1iv14rkYFUrXxOxs7geWhulWhWPR
//5HhkTf3O/5U3VFU+pHPdyz6enfNLCT4NeA0OXX9vZGvqEGlM2C+sVHrW3Jn2KEXnTEUVNQqSuD
dBMJzlvxM+FAeqLPS7VEAXMUGQe1gSlx92rni/iJ/Z7c4HcUaXDpYtq50bOIBAt/GeHNMTY5KPWR
EzfbuRwZEg1f3TSXzXMuzBT3RSdDxNOvdQdBn8nI+CrEoPlb//VTqaxlPdVV97GvoWifMGzV2Fe7
VO335cfuUYsQd4zKNoacuhAiLJFfUm2+hIxNPhCrp21jhBR35IHuyGwMnhyUfFz6wHqOjt28+Axd
L3MBK9cqJ3vtZ1OAZZkW7sIP3ZHUE+y/CVlZ7VRJUDeQEgzhLMq3YrqZlLhLF3Dbu/ST+amP6grc
7Qavk6iA28PdeKRPs6BAn4PkgRoIFf5jJyZQkckBzqgoY0x3oBKvx9YHEIFlfnKakXA5fkVeunXo
KY9IIdrJI6lozKHxys+oY7ecWCj910OCMUhvH+MsaYRdTPZCDk7Ps257WVNM8UTXIDVbtAe3q95w
TTT1ZrgCTMooaQyDi7hHUVPG/0/56eAdcm3PgP30iPyUpu/9SC85AjmBMQ3+GPRHjx6MU1+66Z0B
WaxWb7B/cRK5FcydBjNn5jh9E7PUvF0xTq0DEOmnAIK+u4OmJR3Yh6iKVUD+ySB6Xi6fuUbhrvaD
H01oppS6SrbnELAvp1BFg8yX9+h0WeJOdeFMoSH64gcOK9b0Ohu6jaHdMqywy+UY3lr5Bhm8k08a
Gu8TJVFz+Hb3faJ7yRzjpVu62p1cPret56l8FNsHzb+j7cZ6mKD07YmTZh31UdXQZPkrotGXvwiO
yW7nVE354eO1i5ziCQSufkd/AIEULn7cm/ef6nQM+XoutlmAREl+wHNN8aIrSNl/WUMxye4Ba3uK
RpAmr14fhXvGgEynZ2CAVidcHym6bIVKR4cE5sUuy/v8wFM6BSPgaQGEzWZ1XACNjMK/5Ags1gd7
NCtx4Hx3vi3ZfDyRKy3+xi5QZS9g+qL8cuKN29c7wTDgu60PXLfqP19tz+olLiFI7+wNlG6mXDBO
Y22PjrsaY62abVq7Xn3TQScCX3nXgEyGm/CVoL1Qy3ZUAgIQUAkSeDCq5KRP4nmLXrGGyMytCakL
9Yk3itN0UO27Yswlv432Y2tvtucsP5uJ7g8vw37i5SoL/eFOIIxq8OiRFTqIlQ2UATKXTCNR+cYH
luHwa0dMP8djliyVmwg3VLb9tZ3Bap8Q1RW847ZA9Ok+w2be78enJCQn7gMeR1uzfGGbhkDs7T7z
F7bWWAgyo3JWWGEkrETZOCq7GeNc6e70MSD433i6SFdjG11Mx7Rq308CecbH4CaRPQpEC+ydqm3G
WYa9rA/0XXt+0ls18+Tz9zJVmZvG6GHA9c0rnllN/A+xnpg/O69fBuuIg/R+MixqljKQaZs32DeH
pz5Icq5Lyh246t+9yW2xE+hmfwrpYP0bL7z3K2JhYI6ERTNzDPMn+NRYOiizODhYscspqXbR5fCe
OVibhS1cje8lhVG+RroGzQbaTDv8qKoSUtNGyp2iJxW255sb5KDSXeGLRMVIX8WPkAOrt4Y3DKYj
ib36DF/3EJgQ643hjO82Y1ARbXPfCClJz8WXAlNKROGSiUzcMcyFl3Ini8QilyL2yU2d+u7B5DkU
fzklpOrccnc23C2W+4czkS7x/Du1a2HSg/Qs1JkuE2E0M85Zm2bKC3gxbqzjcRdpUyGm4dJcjucz
l7IF6m5LnD09sn8MQPpSdCk9j9pFJX6s/spXYORU2OyvrFII3OkSjg/WfYhLgKRG0bYsUVgKyObX
5cVctisFBIUt6x4WRAKR0V7CnjHLhUUvIt0PcY7EGCGuzL4GkQUuksZWdYdg1MwMU/5Pk4ksnBAY
Ay/gGz+m0/P2uGiclvinKIHxH1SmJGe1fKzWuhK0CzUgDqZ3bbbtYGcZDH+GpH3TsJ5XRnJAfFyi
dMVzkJsBS0k0YoufrAm9zdYlLQRcVi/1ixLDIqjKWiKhCBCYK29DM2lKfQFfopOzAWRKaOmGgHRL
22dmfjTmPw+zyDyvVPdGP7vc6lh/1U8h5H6yndLBb97pucwhMFSDJfD6mD69FkssM/DD8SZHtnR/
RiJ/KH5X2wtPZlrPaIRxMI4h9NJrEAm5PCqhkDHtJyWiqaH+0f+ONb3A8DQZW4SkUecoo9QVkeam
huOxL/o2Uj7qgwbM6E8Y5FGUB3vTf9hUzNODOV5OBoMdnksEY+8dieRwwhZ32OuzAojAAiLTz3nE
NX6qxqorhrtdLBwbp5ZnC50So1Q9Fp7P7aTuvNbWPK+E169mxb3EcEqBABOPOYmRcf8Ngv2LffhB
YzTVy40ZBKAOPFfbuPLOiFC6Sej7CZ2iHg3JkBqshu77YECtz9UAnJaSYx3Z218CmhtiwC6NgfYA
7tS7jWZ624yGBp/QH+h3dVkk2ypCynypiqTW5D/9S17plikDIz7EdwKv/bDNGb17yNZxxziaFMg1
ZyJKwNtDgpeIky2MQoliRfBwf8xvs9vnUzAeJdZNInKr1Gsze5/w3FV3QQrKbBLLQcxLAEYimi8M
e4KajKkAZ9YLoSfGUCEOjff5g36QECoJgjEsx/zqnAkWi8Xc4m7VRiDBzONCqvbaXCPxA1iJftIJ
4HDfPROiEySOSN/n9U8J71s/dtZgmxcT+2OY8XP+C4Ifv+KrZlRxdVs9y6uWOvRc8BPNqQ/666rE
S3kW0HwAQfE1CAR68Bo5/IaasLK3p9BJ4XCOLQ1QDGhpzexg0scshYItqJoDxO8g0xvhmB9Vn6f3
aTfy3dkllf59/oU2wV4IqRJbp/NbuqljFZLU3fDJftXqshXmJkQWYYwTpXXdVYyPvWJl9+amJwHM
6RTbhuTOcaT54TBw0dQ8fx/H/IB58I2xJLxiGw63dJiuj41CN/tOU4uFBUcFzFddpS3lIJQYWeBx
NSh5p9tdKGkINwfjKssEkh1Ca29QhNeUiSgpTOJhjixVdFn99FdnAAJmYZqP/6nb2CMswD+9PGDq
4UcFhvgDnW8IoKHGHQPArTeJtdu0/QAEqL0l7GmnOGjQjxeVogg1L8aU7RcBmH3zguPGMCWgoogY
ZXGqJUwZh2oBMrvVH1dK4RL5dVS1WmE9VqFcm0NcGIR2VZ5ZN/98gugU9wCdVHLGV6GQGooQcppo
tDNP9RQ50UydU4Cl01B9WAsSpH9VJ2ttvN9++Bnl7I/N4HwTqU86Mo9bogjewVWoq11MUomj7Ucg
BrsChrGC16twpXOwVNRT+wNAxIMvFUUdVoLSLqcjwSHaNxqvNMSDYWdPAi/TsJxdii57JKSyEdIj
2MDhUbkgDTX2CtP0YdH5JAgSmqPF43GYLcLTqhPAQ0LLJE12nRzsVx59tGdgg7fEhoMnO4rEii1F
Z9bq7NoOzb3NpSgfYPvYjsqOggBKV+65PwZYIH4+HFCtyJfmMnZpkIMNY1RKRy40R+zFpiS7G04J
8e4kVYbLmiqi+PnBU0n+JebSKE5Z7wnDDmf1MY4mqPHpmqtqrXR2ubRMBoR9mXnTxLWAMAg0zi8P
rYPe9dxGqO9Zsj6HVBfP/5fWUTVfh0DLL93OaWm3JUggrS7zG5doA+/SNYiYDAM1HwpZuUFMjKZW
ZFiZsIIGrS3PtTwnGCtIzv4AYlf7m4vk4sntTSdB5ZlpSkPYamziICoL5qMXLyabzRirCGpbnKi3
4OF4rb90tiikCJEyp2H9Qzqt5xqjMG7qy2pwhnJgjgC67zY60RtJmD0mPzrcOp8XxdbudZtukiLC
HXrsVJUrZJ/WA0cvlrRSrpKOuXvWgOVoCKopMVTQZh12grLZ22sMs22TlCQlK5eeV+pTYNme5Atd
L3JAaYGRyLTrO/MJqAx9uowqwp2B3chu1ZxToaj2XAg55Q05/MHfYR5BwtjR+OpkPvmCZYYC62ZJ
sVRJnOewDtpqfE4NIoVym3hAo+xzhYtKZLuqIRNKxCKE0ybqPxFKejLHWkuwax87Vl7DAsXfh9yE
2uTT8OiJHNLqVHwVuAduSRX9q1NQqmXzwnlPPD5+MBDm7/6DcVAthGgpnPcXueq8Nea3blH2AP6/
eFLGz8NCbCjApNnkLy4vgmgrz2wFPnXHuxWOPJXM83IMNgUeZX/hYnAevikTOimpPXW4sJm4wxdS
To/4Yqh9XmhQ4w68B1H3jNIuAvNcv7bT68Ws5gZCxM3bai96RYzG7wWNNgNgGz156ipnCbw3qB6n
t+zU3nDNmoJzSjd0rF01ULNlFkX2vO4QvyivtMuGWtHQUH5DC1ow1kx6MGwErmo28sNI3rykbST9
XloKn5IrwYYG1x4/6XMKHS1NT/I2aiamOKmOHXnoHv+7dpYfyfaWdUw3ncxuX7jGwCatsHGkIrAK
E6BNbec83yfFwDAzCex4pR6z8Uw2WU0N0NbjWf+R928iWY4sVAl6e0kQAEj7mqX2Fh356F/QBVK5
JZwqh4J6avvjge6QxCfuPohj2bx713EPzjQIS6QtbaaAoIIEOk988H6OiLihOp0Ze7WFVDwySb7A
Eil6VsqzDPJ7iqVn/cYI4r1fggNU4zR7YMbMQQO4itfvlFDux8YNOsRxa+hM6XEwdmIAZvtsj8r8
+WRAuSrons96iXoQUABTWSBEDdA3tznOLTdsIayxE98wJS2D55/fPWBwxaoWp/lKbYcMAxtUHOT1
fKb3zeyyUqnhazS8IO9PzWkHHZ8aWfu6tjcHUy7wt/O9ChtZoCXqi4EkQtsbuSRtRS8iJdF5DckN
JYMRxVu9PUsQ1xF/JNuxl3ZD3fXe9msc8BEOm4hrND2YLiJzOnoR6iuycNxFlfmCA5sf+j7xYQrO
gJUPe1h0kbpywMieKVV6yX6UEaeB5XJdZD2UiP90S0V3abcUhjEAigdfAHHZ6u4CWtTXdzt69rAf
yF4g1YlATkYl4bPN23JuJmFSQMtL0KaDTgVdL2EjAz3SioJXudDruEjJ7oQ5Sq5FnlNwNhoSw0Gl
Sd8PMjEmSBaAFcEcFerSShpc0VVr4lTlmLd2SaR4PMa9Lx2+Vio9eTj6apE3mZqqBYCQ3VK0OSPM
Na21J9GuMIk5Nq6+DZn+VxFxHlipKp86d1W0EpJzTnuwIDcM1mRzNLm2o0IWqdHLzJKY++eEsmtK
jHhNSFqvhMOlWV9N4o8aeyadi+wVIufEn6HK01UvipwiADqSA5CNBFYzeBuBxVjMTk9MAye3rbVJ
qWqQmqsA5DJTRQP6I8pRw910EiA1Ocztpeks+Vx2u4gBevDBjgY3Jv9nOlfiQe6902IDms5AzQ06
sQjFPTj1ixGaM0rzxZyz2btpoSTBKzgsGwMpIO3vRupIYF6+iRpea3qlCJ6ltKD1MSpsTS+W0ww1
bvaSHu24JqTVMfKeWJ+/f8W+X5BA7+SJKrc8vuffsQ0YXRXtxweRoGW+0DPSW91nXPRcE8NKlZkE
UenTUXT1rz/cZzXx80+hsLM6H0QwXJK4Ae4QjZNjUFE4VblI+yWoJZG1JbQECPYDg6zqbkiiDW7n
fUV7ZhvIaovmbSxUQ60ME5IO7xydZ9JD3nXxEWFZ4SjhVfTcccE7GoClhtCDzuebAsVhrtHQci7n
2WmG4n2j9F/178hlm06cK/R1oFnha+8btgTyhJGxEpIB9Gw2lLQK59wLan1HXAJMhpFGWD4JpfKk
s6gQOsR4RtLAIgC/fIc9N2I46ftj0rWcUs0QDMTrBta0In110xA9XEQNx8nDCsLdQHsDLlK+zurp
qDXgdVxrnjdbdH5OFtzbZVGaGZScPHCONcObb0vo5TdhTKFfeQ6GIuWKqHZG36GiyAZSbeJE2Byj
0FGXB/kmfsf5A6gSDgQ0vCVKvPowoKuJMY+xaDD5V8sjT4Sn4x7jio3W5gUmCkz0ZThuKj2AgFcD
OKaj+17JdA5UmApBELB6HJaQ/GgVvoC6+CyIpslMKD2uOa0GlDHNBu043kdoZcon2fq9UhwuWZ7o
vzPQ7ww8WtbDF1rlZtIe6TkdKmL2l8mPmrQBsbtHB3RjdidrsS/l01ciHghNS8OxcS3NNfhxpPm8
ZB8DG5CkZBgKWSBLtMEXxAOQjcefFi/DL6N2qUnIW64zcmORUGCnF2QcbMd/Tx036oYXWKHljNSx
DokRKfzQV5TRsOksjIUAIFymQtnvw/ASH6sWtjPkAX8VTtTcr4hRBNNFVQ2sn7ys7ekNHAm7JpFP
Y1l0RLBoj2Mw1rvV46vimW5q63nXkwX3uhAkZWRQeaJItyzIglNBhS09WH9ChyROotSDJZrLzpJY
95dZpwTYcc/Qt8jmLwbfrsn2DTMFvnaMDZC1FY65xMtfv5EyfWn0ITdTSxdqcgvsuqynZTY5vIrp
MLl2ZZiQwQnmDuNr+VxMuQVa7MfXIChLSAqMXaxDo1SSYW6856xZLCMyIfWSKIqlepzLoEHvu0nf
5moqv5l69Bgieq2EE5iEICwxEmTR0USqiDcocAJH6lu2g3aObkbPBsijRgalE3IqborKNRNs4nz6
3UQYSZ2wJmrmrJHZ+nfRWJh0lujf8M/kOxvkRcEr3xLQgYIl8iUls0XpADtIlwW246P7IOk8DHaZ
TsMwAQIXHB9Ps/P/l36R4pWj8UbnuW5D2Zx+IodWsPJEAhILPGuVTo0elP2CDHnRuGno68JiJzbi
KI61MFpWjapDbnIorFBAsvoLt9NDQ0tf+s7Am/fqKG+AoxAzq+wCswL3HA007cCh0c7jjPzGiGxQ
n1h3aWqtSc/rzWvXZoxMGuuzl51suMKtwrNZRA+y5LbbTcH/I2iQg6PFlNYJ75r1p40R+1VSYnlM
xE2x9CwW9t6JUmI5kGfEJUK+s1kNbEecay8mDWG7acs3a8udqisRNrGTQjdo3hnW4yOJXdC/7tz3
Y+V/ggtNo6r5t7A2Vk4890Y696ZEcWQtQQOkD2TL6+Y0uTycVzNQYuXOu+mgKzu+p3xtUO8tBarb
cBIeRQwkZN4py9ElECS3PW/2DG1ZDYL9ez3Q8AL8tyih2fU2Esp2ip22VPSofyZhYJ2/emBTuW3c
6tmejl+7ef0a8X+sntOXd6p+PoyOTIhGOt6MvzjMSpiFviftOd4feZiGnE2Cg99/dxOfSWUkOiEm
x2FHM2J7qodtri7WUxe7SgyrQalGWDPcrL4uyHx+4AVue6/kzW4nXOMyVESXdtKlPOGjDBqmkofJ
40aj3FPhTzDo+C5pvMf/JKFJqb/qJ8Nbaz3LUsg1HCJ3NajwSG9FEQICi7f2GnRSUpiwvFij6qW5
PHnoqlrELXftiaZc5cbVQedrOtm8Cq9jUBtDfqcpz3WvZ4WypakmS7x3V9769MQEqNvsopE4V3L1
7k6miUnmKejQNp83t7M7/61m0GWOewlgfg4aEtELJ5I1r7/8uGndBlw2SoYdJjnk4vjIn/poLZ4F
yJ1VAFSwrLqZ8dXhvJ2fTQFhDIXZmkH7R+VDwchTQxH+RrEIt13PBsi0zbMBWiek71U+nV7OtN1W
NEWMSPMdo9yYXwv3Zs5PNETwyrrxylwrqx1jH6GT1WVXherPE66c7SxseSnhameb1ggVBiFheKHq
dWxRoGvEsH43POGLh3gUNVkOs0DIKTF2pUcNUDZ3TdQ70qvwpBH6KCIN4MDquXazNYA7yFZUyBu4
9Cjiu97iK4qCkdsQNmMStQW9+0eCe7BLkUv23cin2/s317i/57W8QXHcv1Nwx0cR99csMx1KVcur
f9MHAEJi5+QmS7X6rPDZVUt7DTDwJUa5Ef+QULeDQia9YKc7lPL1UPU7YI3OgD/Sd444FcSLA7ct
kOnp35abCe+scDG0COR6PtLz85igCJfM63su9aAOaUwIOD6TgKuWxcKyoSm/FHw3l0G42eRnoo15
NCCRg/1K36w5E2jU/jULreR6tlAt3MEOeS7bcxufd1Nt/FUb4Eyr6YmysXYkVz0SmcgiDiQ12ffs
vsehgR+PWKTR86+EgIKmyqpvT8nulDjW44bvL8iqvpp5sZuKVOk4qfbnQKEbAxbAlQ3vDhs8Wx5o
7enzsijCjdGxrQq1agifSUEiFqnhI/rrA8NxC4sPi19fcZrF7Y9V9qqR77xC6mAUD19PBQfMVmka
zj4+4mNucYdT6Zos5HNJAbqiveci6VoDbtB1hJ4Rd8v2WX895GnSLfndFV7ij4RQoX/PIcsVirfX
WTKFvSsKhk0GXtH6IKGTLEJyW1yWioCNt/BWRBB87H9pP3PI4Cp8035YY/jd08wubATWV1EWsj03
EmCmF7WHQA6RP+Jrvf0QLQTt1zYMZtTRhQrMXj7fRD36ypDUtc0Th0zw+HEqmKNvwYwGcKOgceZG
N24wcKWeqdNRHv4ncArQ7LdyxZ7vMA/QqzwftVUpMfVmR2lqXn7eMjc/3oq9JtbkvQT+dKa/axkU
rpPbK9tymLILbliuoLrObXGIS4XXQbUIhOzEd9P4h7dYFZvfjNC1j7ERTtXGbn4avIYkJ8buiHBh
gQ5/g4NaGZ6BUl9vdYfDxjwB7XPGG1wz+Wj1UBMRYWG51JgOb/wB+38rF70Hayo4ulQgU7pEsflI
vruevxEakFLOAooxqJrs1qEdcr8YCbraICZq4DXJA8le0i3+EjLCflrUU4Uyr9Pjear8isrO3gqH
s/6CqNrpI1bpq9Ywx8teUTq80k7l/Sni8Is276Htb1UljrsNhFKqpsOgn9fUKplf2JTRn2L2Tfon
5miVpwjmBUy2ng9j31ltPmRdVSFqcfr4ICZK7Q4B/curpUdxKqlB8yAB/mTJGLmPLF6Mbc4JfSZ4
LlVdjp6LVxbYxqrMte1H25C5bV73i/PwFTLD8kwoFf9qVCkgMygN5TdCXEFyr6BWgF9Q/GvVnBLH
Q5kSwEpUH+uT+HWoIr2N00dGv5m5JLuBq1qE+JjZQ+c9VsTf7S4gzeHVCF91IXlz26RBpLtDw9pI
prPLCueCR1NK9FPwOarI/iT+BWOPsY5ZTP+qaqtqpgc2bZ63QZskw5qhNJ1BX+4UG+p8kXmSL4fB
xP0U0osMaK9lNNW0S+IVu1ZdkHNXaMNgIfyGB+8SqQ==
`protect end_protected
