`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
P/CnevYI+VfqqhsQX+nPmKBbWn4gnOm/GImTZtmHd0bcuumy+0MoBJcuDmby/CrVpPqPozpwjBv7
64p4T+yQwQ==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
i72He7ppLKqP4JZ5LvahVGLV8V98MAk6dhBPSVCsT6IH3Mp+hH/RehiKn5vNSAUXnE+33Hi+kqgS
hOmitlNBqpxa5WtZoqlCAoquuFx+PxnI9EsrGHNN204pRUN6iSBFIVtzqCcv9YSMUtU/uYmlPOih
UtZpLrz9n2760RdP5Fs=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rD8MUm8p/0RoDpxgDfdsDdzKYzmU1dBahq6hbFJcLwTjm7x8dQRtVNmbgxEhKVk3DUGeUpbIFkMT
Meb+Zao8tz1fmARL6/eEinUb+KCw4QuxKOOr2A7FkgInafF0Y8glI8u6m+IPZSpkqwtKshNPQ7ba
BNcQQU7/cCFGv+s0wW1+c/jAST1Lh1HCfww71MbIMbQMnOibd7LRcI/U0GBdIZIpDOmfkF7KIK2e
q0kWcEMJoBHaV+EasuWun946HIdC3PIxJHaxqVC8GUah6MTItWTiW8qQlE5HkINTAx7Zs5I7X0N5
0sL8/DIREFYUYa61YJkMSP7gJmV+Gl2CIWxd2A==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rVkWsdhOW+FngGd9mX62S26qz7BFguHCNTzt2X8uT3ohuCO93WL07BEp1+yO50Yz8Dg6Qau5rybX
2jiAPpl/6qxcSARC2Snyaf2091XPg1LJAonEv4WQ4i++7Alg726IbP+vh89gWHj5XWSp4M/aWe8Z
seRjaatA840d6Pii93O43quPiUlBGaRzip8TCNio74MvKL+LTu0DbHbRbw4qrzW/LiIrYq5k+qPy
+F0l4xBdJ8kSVEF/VHXGgC1yRQT8rS766cW6Jlb3EAd8m9DF5lkufSqdq7nWqc6kRnLIj3/ibgmY
b23u+PinI/PAzPvqb8RJ/j8Afid1GZo1giYstA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JcZPp1UoCCrt4yA2WvlR6PkvTsot25ABKOqtmqY/0loEUOgdYCSpVkXAU+alxUd6otKcmXCf2HAg
7rJPauKXgB+dOneewLpjuEKiNfEHAs3ejVPSCzpE8/JtY8fvEeoJ5d2drJeLhLcY9Jinnrjl8b81
P5FDU92TT7ohTB2IgtP7Zh0ND8bXvtuv3/vC9CnKOizNv+kxe7Z7LzVCaiV1oA7wc4L5I/2Dh16J
PTzDsNDDj91njaZzr+TvqdUFY1JyYiRwq4hXnkkSUugj1sPlKMCjGMOHvkf3+sLMR3nciJ/Gn8Ya
1elaivRmNYwE8pZeeVCvHjNBxZi940kQMnnJmw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ga4hq6xCnjVtTqqrHYBJvIwnj2xO8dzLywvF4L06GkZbXI8iTGIfTKrLdwnu6MFEEfLNpo8GDtj3
9g7sRk0PrGrOjkSzOVFCr+BCsYFN0zw6U0RzndLMe44do7d0Jnd5LFQIwYf//sVx7QwwvPme39tb
hb2cQeHlRiTkssYTTdI=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
i2m2QmCbhCjFBPNS9rfu1JX+Ipu0pZjaBOZh28EJ8U9CudDAbpZhg/c/MmwpJVzH+46PsC+hzkKp
PYIqIwz3vFOdQTzFSdz1SlF/z2+AmlwUoie2G+SBi9O+aXRA+AHb7euo5MlJImVhzbTBsVZ70ZPW
ytwUEzIHGGDDQDLdkXhUSN29YHYcKYtS2JoeqGbkj1GamvEWKkssZiZm0W+7Wag/GqMnleCi2B8H
qGyjqSGiTHyxTZAL7HeB5LzowGg2DrlzBiriloFRWiHd9phKlrI5WXmwkJehmDm2fm5LPuqcrMTn
O0UmW9ij2ZOD13+FeMtYx7c4SAOtr15Ot6XMZQ==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TsDaQ+n0DYr0uZH++s2mUqdNDegca0Md4IyvEVTCRSQ/vA9vBx94wuhciiZwuR5BWBuPXMBvRzZM
QU0eoovdqhm3JM9S5Mrri+QKfUOXVawQvsaQi7NvABbxVONVZfoqqRKNpQK7jcs5fc88bCJqhz/4
n/R0amkr0j0qbilkVTdF7wZHzkkj1qn2yjHoVX43TxPvHUgaZg2Lo9RRitWosGZ9QwQBuT+KXhtf
jF1szWgP68pqy/KLDlpekE59WPd9u3IyMealE8hi8NnsCd6jXKj5pbiVyA9FEHcoVwvHTGcjfsfg
z899Pr1YbXEItcramTfGEODIQnHcPYYsyevX0A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26688)
`protect data_block
jQRgxtBSFDijThDBaRDNqbpWWPc4G4//ACPplttCYjmqPh5s0SVE70mAhlfDm1aqHIwmBasgUVRf
CpTip2INk4nOcCvBaOF0+Rwe2/X40f20iQbckMOqUtP62HIhSD+0oX6YyL2Whl9BzDGKaYg5VZJl
/oYVdrF9a/pcOxuqwB5eMdO2fNccuKWEOMPA/AJDS8QuzfWPXAvjFFEwbMYeloGoDw1Ie6EaD7MU
/C8j2/s7uYmsdGMInAG14MvQ5UyNN2UwP/VzELPf18RJ4jCrnHjxy1UEsPwiwJUxt0rZ5Hx1ifwU
n9NqKBO1yo8h6I8fkjDgOsioD+I2iPXEWz4zXVpErsZbNme9Q4wxB3V1vqTJ8gy9p49UXtymEPz3
elacHytPo+2iqgIbhBwPWJIFbr1MSKHT4I8ZIQE9DImC+M4+GC9coVUekfaRmAEhIC4FQq6p32Vb
sDT5CFU+j1Kvz+bGnyRxMK7ZE20EerhJmdKddVoCLEeJvFjlWcjCsDZxeQmjVpaeQG30schCG3A+
MydJ3mHuND31YrkHWiPzpq8RHVISACGalHWQqNw2p4nlqYTovjf4ubXNLRViaOh86YHQUIcXJk5X
Kp3t8ZOt+KEv0Q2F07pdMAbW6HV9QeBWkBWCgo/IYGF1eGuhp4DSqck/PafupR+yaAn5RY1btJPk
Ne/8xne/WSWkb7WIYqnI4vJ+cqYB86EJYhqCvNSmjCRCZI2fsvZ3TLuoYn7mLdeOmvZE310F2zNV
J53zwHjcw/PZQq3hrFvkp/B50EhNj9XrGgFlp1Up+RiWEBoWXUBLza3dIvb1UCTOLIYcDViybujp
uXA8LXft/D1UoaSheuSkm3uWI0UhFzd2SPlhPRYCIoVLQNrN1c4bq4JBMVyXDkhFsZKssx92c+rg
45PnDLs+LC1b0X6GwsR/T1EI0Tbda0n//vqI+qOHiIMj1F/YcaQtiAVSXr9jfWwYIgkfgYma8FTu
iW9RSumpeZh10WpiudAG8634B4f6oIrzarG+Ql8K13XnTc2dajMRz+A10w9DKTHiWq1G1s8AANfk
ftPbmf87U9+rVx16mQQKgy8IXqeyKsR0g2NVnghd6Hj+niLIag+DKbeCMoyebAWe8XY0Jw9LBJCh
kIfG6fqFUYg5UH/VsKh+Kz3bpNJl3H44KZ+tFkif4sZ+jf65U5Mx0aMMxtDXNl6pUbXkIiCQtWeU
lJQvOMM2ESzi+dydg0y2/5oDCfmB8Sm2SjUsTK/xFWPB2XlcLVpo2noJ/aTx3O5MYfdfTQPFNQrO
f+dsA8W5dPDyMSaYmi+ZJ80BYL7AoAzCVhbCF0g25c+lC4xmOizH8Z1tgX85zil7lyaiDNWBXEAw
2Wa/hbmYjShHK63AoDGGptekLdYxPH4I4mNnKvKUHjWQCtk53JUkMQ9GPIJyuGVoigQc28K3O6RK
t/qoWsR+eeDnAF93TONUokpNqxEsuW4XzPi0UlFFkuQ6vItTISEmu/1z8bZrspU7soI2VUO3ikVt
BfnaVkTjwZnY3BHiuE8EUSuoxHkF+3/prrq2svwUpUObfK+cM9HjZGrC9hCPktg5vL22QY3IRADA
6dDKggvJJ6WjX4IXe2ZVAc+fWMe9uBMhhZ2Rb1p5YCi4gUTXJDPAi4T7E9nG6M+g/zKJPxCuhoZF
sRL37Z4OSxAksS/nRgWMIyKyFCl2m4PAxpayIz7rOnlhjGkau4WxDCVb0WWRLvKihrgm2qOmTGiW
PrDhOa6b31R6mUCDi+Si8rLBlI2ixz3JqwwO8lUgPPcsvdkPflU4ujdh2HlkBEeCy8pTJqtzK+oP
ZZSpMxfv4cj4qiNtiON3CNop79oFo5bHwOwEzylpEfsuW8S49yNvCoNsrTZxj9whoyVs2Yz3CrZr
v5UZhSOpfgyedxiD77f8+eVEspfuw7OBhQXoUYdCO19Dz/DhWg6T5PfaJzY7XycemmZk3r4ar1YM
GqYplrXwr63dS8XtTWLwMPznzY/XY7F5p8iSw/tGYTS+VcFGUcW1OPENUezeOe2lIQpSOquOdIOE
Y7nms8jo9Qu404h8/KOFbvyTKvCnBjtr15ib9vAV6roLzvdQwJqhEo1ZFMx72QT/m1MhxDTaCZE0
Qf2Nn3Qal4WCyZCCvk7J5+D96QNsvk+v3/Z+8e9KunmAbu3z5DF6+qBKuDaQMRPSEbWz76rC/YmU
kIher/a5pspPkrqEeq3rq/Ui4sbQ0czgWvEKYIE9BOqz1VoJVKtDtT+ArchrfiHEtckEJhJ4y1SL
MIGQYv5yGIdOMoYSXfMPyQVhI++LZthDYEOVRG2qVrgFX3bcfd33CdSYVpIgd0PZrBpX6Tsg0YWa
u5rOtNvrNJq7WktCWOwFidtVY+Z0zyDzekCDI2tEJlm73ZLcLv+TGyxtHDXlr5qvQp5LE7WySTdr
DiYYjYMpaCBQfH9yIwRLgEis640ne4iclpnkdVyGcv1c6ysDZTjxDFRJkJabUxe8E/Des9HX9GEN
Jd8GbgYNPE3SfEDjhcDDed77QmT82OMRUGLGLrrFCXBWyGk7Abi7yu2AH52GHBqFAZvYhGXjNw2i
gKzY17LPTU/ZFRQ3aKaWY/gYLYMFpQ8XEwcFEU9jI+6RaSITuu90hJo1dr1ozz9B+ghXinbvDI4j
1vViCLO8Q4Znl3YKFJqUi42FTGfp8s6iqbO8vfmb45J+CyqCVEPnI4iaxYBe6SWDXRc653/jcLn+
xoK+fxG1eMYZHAnfzHh4FIPRgYvn+tI0Q0V1AeVVo4kvZE2s72LwSmePL1nO5K0riZ7za95X/Ils
aqnvlbv0kplBEjQjXT7EZ79SvR+djQLxXZfhXYYPmtCUBbsub9ow0Y0SfXUMpXFPuYyyoByq8e/Y
lwz6VlgLO15zHAXtOTtRw+7Z9VSyJGo8U0MT5YPTF9bCLaPMuHNwGAFqVBCTZlW0l1SI6Vw+VYAO
EkLNsdsEdlxHyK56xnb8sE1St1BkwHqE+nP69a6lmMgHd1thDQx3IXbRaGjt+7EzBFa6OXaP5pKf
VUDP2LpxfHzUbS4FjfC8fEVBrUONioi/uOC6ekaRGfZuLvp2BpeyRQlZKo2HkELqTtSLY7EnFXMc
m8hC7DZW50Pu4PL5XpZ/Mk3kwXnbVGG7OwhkA79fbulcTvygxYJhkzDlxsEFe75EjGC4okHsvf/O
qcToHlVsSaXl+oMHxsmg3kehITimdMF5GAicn4O0AmABY6l0RZEhRmz/MzE2toSL011l8Ka+GAsO
RXH0YAY7GnvBpxfymd7cOSLKYdnXLPYrQrW+AMDtl5qfG22mJGudRJy4sKcO0PVwA5YeOZpV8ckv
at0I/n5I+EOJHqt/9SvwALG9MbgJETFndTILSP5SYtRJ1OgoDyg5vZs7Ikh2wDVNhv2Qbz58WjsF
KWEOlSp3z6bErZBK7kzraKWNcCM7NUlEkR8SSLB/n8ZgVA/BpD93nUKrdFWDgA6ejPLm3qK0yMzn
ARYWzhQfpevfvxWfMSSoi9qJETdI3Ta9QKta44vRQF5q7/3S4eziTptZFxUYewu/YDsWpu3x64LX
AezUu2Y9HXG+OrHRz9seVURznxA/+37p+zX/JwmWZtouMwuBL5sljEwSkfJzkZuUgQUPjJgq/2wL
1ZwvEbcqYd8XOxL2Bw3ZiPuRNP4Opn2uf8q7L6o61Qe2w9MKGDJ0JriQ6OPucsNLbeuotEJnlyGa
I27anyF3mSFXdA76BgvbfKiP/M/DoCaCjq5xNT3l/6koxa4FWAhvAsdbw5KsHMQuNIb0sJkWF0XG
PxzV/FQkRBJ9MsAn/PawR7KWQMLWK4wggi1rjosmRgTrH5+UaPMYMyJ4FZoGsjTIv14fkQwR2+O5
rr+yf+sD3RPesbW+Z2Fj4ujczTeKcNa23uTaeW54VSxrboOfl76BaJxcBVRfg8PgVsKIKfk4q521
vTiZ5HYDljK09GlA6fDHO277Dwfm9LWwjbQHzzcXKqvtb7V5IbdB8e8H4ExqYn+qSKLKbrbss0fv
rSv/3feJvkGK2l8+X5WD8cmkAwFygPkndc5RsqD3PgOp97vXPFZEfTRvemLFKc+vyeabmKpnD+t7
jJZVcY9XSsbBaHHb/vXtwDlzCc0CX5IeUSVhQY5TAKFPV0YP3SzPtWAJ3o14O7TYridVdkREQJvk
tjp84EkmDEc5FwANAvMlU7aygwew7jDvTZE0o7ywFKzbDAzsDKAXgJmChJsCnX9euCR28sYwMoMB
yQDsT1GE7pczH+Lriv7BDvzrwpmIcuQ2VliKVujILPXj6INLYZuSb0f19gnGjFejE6Itrxm5F1us
jTK9nX554dakj7dFlBfZcr0jjRvx2wdyLUUngurc6UvNSPGvGohKTfIESgXYJ2oSPt/Pw2APGlXR
jOxr8wzcq8An93VDDpf8bcjejvkzYZsvkBvL5fWcPG21zKoXbFrv+uCzWBS7Ww59Zbw9kmfFMmcq
JE7XQ0gXQ7deAudJF8sXi06A+0N+iOvy5SA7eHI54uaB+Uax+M39fDKCPOaLKp7sx71Yg3GxNozA
t669shJgshDxhQisLRKw9Jfj0eVdI48WS+jZp3u79HI+LmdZNGjyIjFnOVqFCz/hX2HHLtOnEEtB
4wSTyxDJXerwfEGUEi7XMHIP9VI4LOyIbNa7VIyPxkY3hl+h0Xqzo4e2iQWd0FUzAvRDmlGABzda
RVHOtKe/ZJPv5r3ff5T4l7UbwukgpFRbwfsg/mHSU/vhIuI8RKl8bLwIC8LaJtrAyVI+RGOPluX7
xn4Q85RPjWr9i1rglDuewqCgZrV4P0lE6mdj9JH0XV28375zOBO+T5IW3O33BrK5zXLAkabE1m4N
4/LydsLsbWRKy0geTOdDWNsCbg7hsXGI9PpFgyptr0GjuMPdhapO4f9/ZDfgSTzMQMsBGT31iJ/v
GeWKjUFzunvrdi8rT+vqWLcv5B+ZvpD78dzOJQGx7W60Wwf9ASICA4xxAlJKhKZQTRFkub6cUorl
nQNcvaXsswNQGqpwG9cODitKYWBDP4m61a5+etIpLuIpCZEfQqym57/MsrefisDBttDiEhZVr8RY
i84ohLC0SD4bjk3E1sXzTYmjtUbCG2VFJn6u1jViYbj3n6YiyPA3tw82R9KOiAOzEaii11yJfzI7
R4MTnn4FKznYRIOpDg6+RC9lZj0/mdhQvAyqoI80xfTdrPKFFBS8zbslWSRFGKgrVR60wLu9OlZ+
aMNP0T6uOM8use43IE4/JQOAtio5TDmcnEbde/l7/3YWL0FQWayHA9Fyk2GQWdpOwchEloYldZgb
PZubT5VuNn7pxAqLddoR/dgGJaNh201a+rQCRmUIMGxkdpA6rjPVNVPoLvmRtw0AMfGgN/T2GfYX
7sduDnybbhsHdXesDfmuHy/FGG/oHcaOLlHf6DaJc4JYfK75j1NKXVZzPtt1olBYPGW59+h6UH1V
e3LWpIGIHfNSFnKi1/lpbLyy06hRWVd2kEd8/FhlQ3mLk+whe3wMku2+F9ROz+HJE4fVWNtuFNai
3Nq7n/nQm8Lsec7UFCVQkUM977/TSg4Yn6grZg1mcXv53iMIxOGHlSFzwJeOPDwGwTx40y0GRbh+
aA5QVQ0gnVz8tLb4T7KFCWSYkl2PHMyk1MY9/cUwG8em5GhErZPfNx7RdHN/T6eEUMAXpDo/cB50
D3pMxYBUadfQ7tAzdQLyekMOWrDGZccyObaX5ZpprZ1TibCpLR4MdKwZsoHN9Ku4A7pwsEPhsUvN
IRXicjkclWaW9YOYZJL6Y1VVAFyuxABO67Vv0vHJwtmN4itjvCNUAuwrLy/7eRLhV8w5kd3S05BP
EkSlnovz0ruuJn8JZAx3bm8lNXs1FMHXv0cWdnCSHprfv5dNEtTcGD1t+TL40YGfZsBV1i+HMvA7
VpsGbBB0aaSrMfWWLkZFOzl+h6VV10WFwizIrMCqINCmb3kcr1b8ITOMJbTDZDZheKkEqK6prOPQ
2P0b7HVFQDPoJUQEkmPWQownOvW/l4zLouOcyKwhm0Gn0d+WzAEJRDMCnUhExaZl2RK0IXD60r+P
ofPqr7ObasAS4VHtE74X+9prh5PwmSZh4po2PlwbffejwmLgobb6uTQx7VuQagu3YxOvi5rfX1hY
3BL74iftLRC9OklYtk+KLwIqXgX6cGdrSxfdRuUWHQfrSk2jaomrgwwKUj4z697vLmTAd2G9wN8c
kYqpnDTbUtaDuihOJRmZvnyMgoG5pXn1z7xxky4Jg+mo2z58cB80qnEFidNF79OjPmMUZ8jQr541
uw3afS3t2S23jUnc9etoT12JpCq984QLHjIpEy69zsIVjpP9+2ja8Qzsv/tuIuQ2eoABlDtIO4I2
7VqlOfbv2Eg4AAcO0ubVX7eboDnEDFzhGDjmKyVQjkmLNNy59NIIdeUSH5NAN473aVAS4S3NxT0G
3CeaDsCoFHlH7x6Ca4y/Jh7/7EoVXT7bpnUxHxoA0wtJ//oQ0jc3owNQ6WW/CSF5TER8g5rL+Uke
LZiE97h+Qjd5+sYXNU1anInjYSy+pTvCdUqUDjdS8Z5pppcyQrGQpwbbFNHdf9MX6oNs6yqZ5it4
KUmiYzu9eMAWoH5PLBvGOzDeGPPUpRNMjM/mHOb3/choEyJn5tzEjk+EP7YOMK8CrZ5lOfnZV1mK
1doVaLdSza8CUo93i59Tw9l+lqUL3Hm03OAvgaUpxwrDvf4g1pMCfAci6fhDRrOgt+8XXKveUB6p
vsei1t/SV9jsLfw2L4Or7de4HTBlgyJkjdeagqjuj4wofbixrXEGKa5J2JxY2OFafqswtGXJxW9h
JDilF8arQta9qbu4mMxkuqSiqhW6nkOn6MSzxSEf1NSiNUgCv4W9Jvz14+fRb69qjTifv3r2q+HW
blZaoMu7L0xBc6Aq+F+kGt9ZotTkB6N7ro21QW7MUvxhy6aGgrwFM6FeWzOpYZS6qkncazN1tFJJ
c2YF9mcZT14Sacg1RUIfXKeLh8clpVwG8CZonBLw4H1rI2OmSigN2wpQvgqG4StTJxRkNYOBNnRH
dBvO9J0XRwxxLYCDl/jV6rTbwRnPlCKWnBkp9NRXqrUA8yS5CmjyutOWkmdaTXm9nDNdhOxy4VfJ
O85V/mYZyeKH6gCT/oz7Ork0NF5cV0cSlwCXyep2BPejUvAcwMV/HHR85XCVFp6opmE44jwkxVnV
KBnVlK6L42QMJ1CZXc0CRR2YWiANpYDr+9aK7MK2zo8vO995tALA1tOuwLS0hhzKf/9jkWxXehS4
L/NgbkvRzro1QEYRyyMf1Gt9+LCz2OuJHQsMwHlZVdYs23w8sRcY0LYY38cLMKCMKSVZAfXa/X+f
4uIJZsep50KltAIKRM1pSzb4lxFDhehM1jsvHNTUqst09knCEbWCjbVaTr3wVmYT8g18xwSI5yps
yopnjTI+Ix1/z8pyiCNt8Bj02BtyX1/Ub8ZSKEIsOwe4b3Uj4Lqq6KhUHRZz+khqwHMOkZ8ccJyB
2+H8EvJVbnSt3LXr70gYdCOtV2jYA9YIn+dfizwnPE03z2OFrXl0lvdp28fPf1RRejC7p8z3bGk+
EgLBjvFxe2TBihcww0Df3uASdvES2MOaW+B33LknY9asvsEcSJaG/uxrgyo2lqEJEEmZwE5zMQnl
OI71hVWdrpAVJ3MRLQjW0ebCaWsE/Awmi9exMUlq39qdpPYemhIt3u8RGEC3gJxjlRmfR3o4p6QN
x6Fb2wEYkIzAvYE2PB8l3X87MEAxi+SVmy+o1bLhNCzRtVjZk9CDaLqosEWz9av4ckXRpRTMDPNW
d3Rh3+fUs3ApxyGOf/q8OgDVuwf8RaRhfVQ2RQgCyEKPc9J6OuQdPk/w8/49nbOu4FNAnKPdnYl3
IRd0/1coOUgwXubl+OLngXFO9pNGPhWtVoNTzlujTK8ojA4xbRFiPFU17+lRl1wqUv42PVAXNELe
BTl14uEpOnk+S/u85bGdG74+rUqBOcBvyJNeLJqys+R9xCIVzpadaGJa0Z+Q5nzxtcj4YwrizOu7
MPW+PORXrraCDRwh0EXhK+C7t5JksOic1YE8+dPiqdEGWq32xeySfczpg9F+kUJXAZnbh/5JHeVw
0auiq9sVcEkZVSccEDzXWddAd7mCQrlAMppZRWv81y8N0H55hFwsEiF/lde4li8hLlFOG2gqaZnW
G48b7pyFf+p62D1o7MQRmeYWGdiJ3IE7ixgBc/CrcSDCiCmQE7i33Ca4D2Y+wamL39v1G2mUIPbT
oTNQlRy6hyVt2OMT+eEyjC00gCJ+QHWAjuoCOQEHSf0wcfGPO94Jma6+cWTTFid2DASHWSfR3r2B
AMZLb6kjciPTG00hp5xPWi1hluLXLApZXxUMkIehCMsUISfjjapBz2mPelt0Vujj+hgJ1/vP0SNL
aOZueIjocO0qAwEebsVjfYdG6b5XSpp3L7kiOlrN/T5Bzj+bCLCk+UPbBx8uFjUkDmCEGvV8I6Dc
C7t9T0pojjAq0M7FH9YpeWGM7jIcTCA1uN+kndDbx0lhLOj0Q7OKcbPbGFiLynghWZMfqr+SWJ5s
QKDT87WMykFu+U/LukAS+fVux9rtDFff1J5SZKd/1ZE5eRUyyq8DEoOP5KJoG/HVqk2QeC9kDYRK
0FPdjXYHx/eNmtJOAe8Z2UBrNkwwdS2JdLv6icd1Z4hnm5BNnSGcseEj3qguDijLIlv1h6f6TV8Y
CJDX0iA9JRPwVhJ/RlIblz+H/kAYFtyrsnnjN6UiytCoGlxNNYZ/VMamEiwgZR75/RWn+a/vX0LS
oyfzkA7qDWGJL0jXrTn+MmvUtMzh8N/JWd5pewvFyU2ymXkWHoXJdmPamXkI+PpeoYTIDeyGUYqn
3s4IGevPD7XPlCLrnP5+v+3/+3KOWasYFPFkgSuJIjgz10qC124b8+8oUfJws7bkfodVoGs5vsUs
0Fc7FwWSYV41JxcY8FT2IIufjPrRIdCdvDIiEnQWSYbMXOKDsjUu56t4PnLUIzyh6/b6Wk1ev10b
7AxgmxdU0AIBdki85p4XT3L26MzC8ga1qbghT8GS8gWILZe+YL7ugLse7hBszu9eXk1Um1r08mvE
hgelTVIXJubXigzG701NonXlZfNQw+pNf3wD2NIs03iXQfzYU5DvonnG+fsH+2kHZ3JENaB6r7s6
o8B/t8J1hclRW2kWOFruliVkNKwhpohD6QEtE0V6azLWvneDiO2eStOypd9D3MGWlN/EJlxLRGBF
klKTYuIw0I53ZhuxnunmqsVfgiJYrXE8K+/m7dkGdIhse7LgpEcmQA6DKuR/UlXTGtNlTciLfNYX
hJm/4E1H/sC0J3XrPoahI3wx8qnha0IkYDRmNBG8VszBmrXU57SQ+d+apVzH6gwMWeIIZjPc2ezx
bcPPJTtQHSmI/43WqSGQ7bF5c9A3+Eiyv8KjzmBI/+AXq0e0ZRs+sMH9jfk1cVVkQ9QtD3NrJ0Er
s2bwmB3DQZb22w9JJ+dRLYwjVtZ7BU5pIlh+8ashwZlnFGG7j24im9Ire1I4gwlrEOT9zR0Hs+md
POmGReBfx88iWrnFz4d5J8q+fz8NvGsXKSXtft+WJOnlQWreNBZA2PESlVljZ4Y5e0hgCrlzuzCr
A4B6r5VcypqA9f+21mcv9H39rLmh5VZOWPZ3PbnSA6TANYI0/M/f2ZFjTL21le22cLHB6+9il1jB
JZ0dO8cRkA9sc25ndDWDXtd45mfM74aZdiqwd6j/XpyhitVbMLNfBkRn+FroZ2ajH6CYJM3x2Oaq
822EHTn0KPHRr7i/jtrnl4G0+Ju2SiqVPlH2to1zxZJmmsW0I1d94SWAwBnsPCoqr3171w16s46M
+syrXrXPpV1hGtmduoEnt1h8iboRyZCG20n7gjzrI6asXGNlnUkZ8II32+6g/Ow4rQBMVrBR8j6b
YGLw5WAQCCQSDbnpVP3GfUx+004uTQ4Y17uKC0HlPKrCALM9GxaahhqdMpFAG8sLgKmdY3Pfdc+N
S+34dUlaLE7UORp3dowTTkR8znBTC0/5wvSt0t21WpOrpQTG+GjLaQIJb/FJ2c2HT3f1M7c3roNK
dgmslZo+/qv0dL3pEI90GG8bYfNAHSAKsQgHHnxFMGrWJZ9J995C3t0GSTnqqmUiBWUpn1gna+js
eXaJi30ejLhiNzeyv5L+rB8mOfe5bPumpRnO+x4XIDz803cFowOFO6NWqRvey+OS+9qTfs2yR6vw
ZFbz1kD3O+tBgPBLQ9XgtnLHRBu+AgQEDeYXYONc6JQv1w7DeqjfsPiEU5wMHx43jX2vkIV6R+95
+7EjhRqGnz3O8aDRHaKtcASXtGq2gDwXQIy8MBH3g689sRy5PH4qRLLNDiSgFLtBxDlnNAyYB3tS
wzD68j4NzmrZ09EnYXrP6EibNf6uFQA9QS4n5FKxngU3tQF3TWHNFJynwMowziKzyAV6IReAIIgV
vz5jiI8GQE0vmr5HrpBELqKA4IYgulGRUnyNNHBf/Lg1DaJS/59Qch5ivA52ncVH99CjWLO5aNyB
Ou1fyxHxmBw5thOMAdy1gtZz8mySsRmzQRGHDG32rN7JRHbBva5MWoYu3W5RoQwdI6sLyoCZkiqp
MPGZWDvBJ4cbCqSCxJsU8fBEouM/JQj7iOKM7N9pu5gDCUidOtvyCrr3vNAMLvbsfkz13JEvY0QK
/0pihXZEPk9//5w4NkB3n+LlwmMXumL8N8AmQFn3Y+/Mk39Gbn2DkooqshvnczRFiVVn1hRQB7Hc
sxWGaEg4zNzyFa8fF2iehGUEqM1352lXjAnY4YT6rTYqrHYBuEeCIbXvxCv3SkU1GmPiopIiFlI1
yO0oeqGaIPMQQsqglWWyNA+zHutJo1pw7rcfvnTMnqlnBdfaMTUE+60VGKrMUij20eYEw+Lk7ptq
0gfTUbu5H3Lpa3eteA5oueeHTPDeAstnX0eviZH/miXdDSYfSzvIZ498oBgXWksrxhhU/ghgkqBI
HmpbqrMqZEdeYF1VNYV7nHx/Ia0RlQjuOLj6ofRwNzEUGwZbtW5Yiadzp5W9dL3UsvMiQ+04sv/p
6Y+R/W9Jo8coyEZ6Rw1/esXs4izTQ+aBELh2JVFoBYNCu+ILmtoNeGXmUCJLQg69qSW9HxkFn4Ht
Pp3Wazs9uAb+/yQL18tf+/eOFVshyx3qs2lqq+fJNG8OsTjSVCpBwP52faOgrQI93wWgzXa3M/VE
xDMUvTJGuAGTBa8l6FlOlaiUda1RKjcq4mxKzr4Ql8AOBcOrr2qOZt9rjkFc/jLCHFvwgvXjYC3Y
hriDJVoccYwEpbOikc32v3nx4y5SuTnzEkKcr3G+LAxq4khSsTZMEJ6ph0d01ePlI6BVlYcTkHDY
bEOTCHlZj1nsAI6ruff+/7sSMyJbTy4YOODWvvu2I1FOol+1CyceLOvG4/JMN2aQHZ5+BY0fcbvN
+4buLmHceVBX4sSmZRpRzW28JkjdZ8rxiIuy1JiMU20Tlqvmf2xBE7PpqELOiALJS/0tnkcRtYeU
ilkiKmpQbLG1bQsvWYD9e2t5KB3nynACJt+DBzNI7VISQRilHQ0AaYsW3oeyzgtNX1mjyVZ3WU3L
vDaa9GbKDapwA/QTpcMP3qrjSBtGBnDpPMTo4Buw9jxmY7kTl73cI+dMKa2sg/WV2m5glQkD5n1q
fp/+WEyYfcSyy4b1dQoi0bqBawPbwjF4Anm5/+cYO8mton9fdv+6uHyyCyyJer6iEQajhBMcFzbT
g1d6jafnSmlgvYiCfmeCl2816Fak0Vp7Oh0NpiR1XEEbo0lgqEy0yieKtl3Vw/aL3HI9Lk1JdmmF
kRPMen24+YvRHadRb2B251TtSXaR4Ao0+BHAfMahCzhCLNgFJEfHHjcAqwI0hwmTsBFJsPwo0cRP
LD68JxuJftbDNfKtqmXsvmZ2IhGJ20Y9B63S1wt8A7nAOYW/+KoxiD1W7fAvKl+Acwfa4uaqBM0j
YZii7i18wov139F9oZRPhvtSupnHF16SugrDsolmm1+JM6kF1aCtMwzQRq1ySUibQD7RW0o73Ydn
nfXwjB239JT2Mo6eVrmz5I8EG5uTNA7iZFqFfh8C2zP/eiBYGBNLOSSm55mf8Br1E4bApS3p1S5c
wGJ4bYpiNMB4DKNhpJIx2Ljp9in9ZuZY9nAxsDT7/E8yKE5ya1MHjcJBdIaJAmgKqeCuNVgUl2jZ
elpzLT+AnjAoDT7dMJuh5irYfyBpKQ3DZaTTedkivd+PCo1XAWx0SzFZTupjRo44U3MiiEH4RAKh
2PmhGLelRBvWg0iXlZXkfMazb+e/4bBl2FXmhnHPEU14iHzOOV1ngbfR2gEJ8EN2p0VDjYCS/BfP
2aaQKMsHQYkAjSe4PvmTsGmg/SKR+XhgQr7uCeWLV3BwBeSsklimUIPbhH98OF6yHDWbyQ7N6iA+
Dy4Rz6eYmrCNYi8E06kXo2IGqrC/O5/D7qJSAPrYcA/iE8URp+kCjZTVamQF9ciXN53SpQR0xhw/
3B5RlxRiVrXSsdQx/MDNWoiAtvc+ANfkQDK/1Lk1PVBNoor+WcgQ/hQFAp4z8QrtAgiR7bhiHybD
7Ll+M228O9n5XsaFB0haDWIoxo4zCxldKWWqpqPKw2Glqf6HdmReskMl3xzenAwuQ35qh4kTaRXH
Ocvh+yQjdzQau1Mq9DiM4rXPzXgJg74MfAVz9ClqojOUjRWpptDTbt3mEKbSaIgCXtmhywNqNIh1
C+EIIPQ5Tk+BJJ7Frx1Ig/Bj8DPz7FnESCDw8hfhK52LTk5xGK0EnJ30hUCJV8tVop/5/x2A16qT
lyKel/JK94IdO0cDmF7twmGBCjvk96KXjjcEzwMvK1OWxeEMQueYYBz2uCAF0BILSSydLcGUfHwM
T1ZJbVGczuNt1RWUNXfI/vqWb6d4OTiuwDgnIDpV7joYKRdq+Wa+huwF1bUhYDAg2p1lwlF5PXrY
24rmYCNbmPHirvFxKz7t1wTGhX7iqsNwa2BUJggh5OBnP7GpFFIacV4G7ubZetxMXvilTVI0J2ik
06ojtsQi31OVHHCmpmKKwT0YrEmnm3McRHoteVVFHPNJG3mClCwBpvtHPSyUuw9jBvN0Xs1ybtU7
i6VORNUM9MIoCjyCxhZmbTKHRroSQGrYFFcN2FTNiQVpYb1ckSGdUYjUUkvDsm1XO9Q6/XhYcUoM
CPTDOkJ2Ycb+cyhB9nY4I+7YKcYyKaV3H4Y6OIxRqk46K5hGDA86DkmYRo+VJ0Q1qRYFyPUwUh4f
OMV78HmVJICiChMipRpAHeauJ/pcOxEXgp2Z2s5twIMazBlmMoKTwJT20rJvTtqSKA8GD8qJmeP/
dNgOZT2XMlLogVhHGVMCqAP/o/dfty5IcN+mVVgLKgimJd/a8bowyDDDK55pEtebZRkrU4C+AQHa
FXJLz/F2EhaPtlClOQTbJZosEBeFOHwwc+aHTUTeHMtkKwZiNdQr1pkxSWLMFeJ2a89xlTOeGLFM
ovaTc45DdlBskdbAwTUfW0Z4sjAZA2O0cKwv+OSd6NlUpBMu6orRFghAF0ti3itvkMxsyLaDCHAQ
grTR44YqY0MDuVutF4TR/A/B+uyFqvm53xKpRDhlCu6wlFsN3k0PngtB7NAXTcbFtg9EuiuvhpcU
tXz0B3Ma3moUov7MhC9dCBjVGnnVi4TgaTzv26t78t20NNJgIIRRrJVspExORjdIeD4g49oztO51
m/HbGCa/svErfo3KXy7cSlVKmOd9qrt2U1GdIpbYeDjc404Uy7MeSjoL6noI/JrRUXjFqM4oFZkf
HoSyLT30ba/ZIYttdjnsEe/X6W6htzZ9eQC8zv9acDfjk5eGIAIrrVpp3htIcy4dsDBX8ZCSbMcA
kNuG3oG0WnYt+VsNUnrtbm+UR7q8MRrNtgAXx48N73CKQGQgx+9oKYxjf1rrDD2HU/eaKaTfeCFe
Nl8swegMR1pE5ESVR7maYQFkflhvV5NQjwf1CRs/JxKIhppvJ2envM1N889lLxKzr1ffrC7Dtga7
lNU+PEFRtY6cBcHuz3n+s7eTOEWhKICrThN2ROW+17cbJ09cC/oG8ChBOGYEunb67AGd3nIOi+wV
oJ+RluNxFyLAxQspHajJ64z2Bi9A4ZDlz4mM2VqqOU+boDRns7jd1gGpin5n302Aou6pM92uYau3
WRRlisKB9dIrZvglOW81aIxwgbAko4viqb6Pv3JdJdXuTFuebkdIPT6RcxWqS6JM+ywTWQX9OOe7
vRU5p+MtA8K+aVJj72qK5ELAeG+93h+vu14uyn9/aAxb/G9VTsu2rfcOQ/DajCjvR/Ea5B9Idv90
5jGI4IAXETSMYTC2CZIziifweu1wysvvzOLLXe0o6netjIXnrxj6+t3Jw9cqdYDHBNnx7Fj6V9TU
7R5m1JGZmFm0xHZVBt5L219nCNYQNY7mHAuWgHHIIHGL5427xs4qd8IiFDaAfCNQmLx2RmX9MnNE
OqoWKnKOaFjiCuxUm9QLPFw1PKxGKREquTDAlBA0kzOVPYt3YlTTNNz9toykZ8YjcdTD1vu7Kg9E
yr/WqS5gYOzr/c/dC1L2i2ONczoz2HGjII7E1aGs+rpfDbN2tatPksOnEacYEXOZVBTlkBFTScix
1Nm5MP+oTWVxTUYK9yLm392/MFcFbmz4lzyH3Z+i3ofuJ1iTPogRajmTOWDDpM5jbsAVO2gE1BWR
jr6Y2aKitJIljAU9SkpT4OGgN1euTGT8E561K+QCw0tE7PU0h4XohXV2NuKAfm+0Efve/xjN04Fp
PSx1E9rWrx+5VFVD9oVgaEAGZ39lVRf7JVN3qGTS+pVknhiIOjnmeb/0iiXnjH9KatVkl8Le4o38
pgLRiW8nokHoodYDmLW+pCX51V09HpLM5vQYDXl3mDBLZOQXY5XJml3pgYvos4hoiNU9fjDmchj/
rCppdbvNTrLjHdDxcvzQyZsgBBUZtFhUhnpB5J/aSL7unDUp0r0kCNAtLSKBhuOYCv/4juvyx5jn
NopUfh0o3vXJzqb2HYdyubaz6bFRgT6EgXwYNr8UutHVQGxq+LmONqFl6yzkiZXr1q/12lR38BAr
z39EmEFXWHQ6fMkoDCDD2n5uJN/zSRc1+LMI/fV2lvpz9k5J405DUsGMJ/D3G+5AtLrnp3ZRE+dB
IdbYnaNXA6GfdO14NT5S81Jt+BNtIHlYIhmEroT9ymRzsTCL4mgqC4PJiQvY9a8JqxbOC/USXenh
PA32M3+4lrcoHfE4oz/eiLdc6prgpP+JodU9nN+ARTReGp2UJLw6L+dF/56flXpAYKTNP/g2beEK
IA2K27uvqxFab0/Fi32XM3CnAuRyK09pgM7vwNvWwJO4ycuxVFsEgdo616OKdOqmInRDCzm9nLd7
fPBaB+C8MoBOsLG3sONHx8/abOLQQEiAa/QZH1voV/ZLWfSRch5t+V/dZwB6zEHm5pD4+oV/Kmt3
a7xzCUS6iH0PPpJZHFf3bPX+FzJgs5y7iyOp57OQe/QTp2jZS/wmzo/dzEM8c/t5RsQafygie5vf
jZ4dBtpku2WIQtqYMbHvKwkuX8KkCXt2/16YABNKktSCwXwHYq+1ZpG5EHOVe65UYgNbB4sxMHqC
MSZKIfJd81ElDi6bPOxf4CV4GYESQ3deUEF9A4ODDkiaMFni/cFpl22C2eFtwqEqQIxwrlzMJciR
RCXs4xl8g6DfSDBW9he2FybAAOrje9sD/8Ji8gtHMj3jsqbp29V68QFBFYWc5+h+HXVCFpFqw1L6
6jalWIAgROKj4+HQLFm0ITRd8JUOyppNTok5ZGGhvTZ7ACifKehp6OzhAsB3uYNbzxiyKs4wbs55
suZVEFZ+TVbrqPNTMyZNn0lKZ3Qu5/tNVpYslqFiFUb3JKEVfazn8Z6TOO5hTQRQRxS/1994uxdt
jNeKu0j/dtQmGnCqrneUTeoorjgYaxyEBpamzRzKCjTo3qCXUWimvJHc+D/QgFnt4OJq4CXxYRL8
UvxY58AeaTCCPQtLhQY4edcVPbi4oeZeOcyM3lcwWXWVJ+gWK/kWNddeV2fJZbgi4tYoUOv9fNRI
pvTd7pdwwTfy4iBaDYu0Y6BMap0Xlheiewd/Hnlw+IrE0AmGRLtcxByZ+MPRpMTAzPRiVvhaW202
iYVc40kYHQ1ihqL7zHaYIxDRism8B38k2f880+EpBZCSQAZgX020WrMP0WbVVYYK+xc5/yxC40WB
SXRujxDQqRmnlIRneCXFiEAlhFEuMdu7GnO9fTFenxpu4fE+zau9Sv/6SMR61Tq5rmQANUjt6Uu9
PFWVN5nC6caFcQOddMExvUR6bUWjKCRmPCU5q11hjQ4QXWPIyD0taSR7jxRJPvpd1X5bwHzhl9pZ
db4sBNmmjKRzyeo/iNh9kVRc0sEyXH6kw5PshGVx2z+wGlvPL713wff3m7xU1zfJRPHjkxohnQHC
GYBB24EYyf1LFGrxUwkm/z9CC/Zs94m4SK/ySe21eQ/GLtaBO/y6CD6ZGLta7ET1CjejdIEHQ8ji
sXuvdTDCwp8DxRbN3aqr3NTTyssBI3Xuyi/7hF5fteEI+ox6Xpr/auJqISvejJvCPGYvAtqIdNMI
Qdg7H3oKDbZmKP59UaLeZOhQ5n/2dfGcZ9Tu3ysaTTDy7CPNJIQpw+8ddXI812pa87rcIYGBIjuB
gNqN7HvWUlDeDfiAbTRojw+UYo0jMm6IZMP1oT/8cAvJ8xZoQ/M/UynjUQhosa92IW/7yo47eBkO
QuCWaXR+pB67tsPoh7Pwq8QX1Rg2BCYviWKxFiBN91FNZ2H3QRl5ba+9jVmnpbzVMaQZ7BdbwBqj
0zv3/VAbzvonRKXGevixbZnYRUnaIQZCjJqBbFhvnv0wOGgH3tTICK35rwXIZa6xASJg64ELjsmY
NvYhEkKGFQA9n7ULhRHpXlQPzkfMjv45++jluj57ku16UkVVEfvbDMuO//s9Z1/FsfkqUvtqMtci
ErdOf4HJay8m0F3TutB4SEKQEr7WG7/px2QKSgdFHQXSYHEkaVGNQXpBLeWNw17EEqV3ItXN9jc9
q6A9VhI4uAIYdCynHaZEpdMHW5kswDhsJt2jGn/TphU2gIb2QQ/XCXJPs8FPqmvHiHNMb557TPw+
FPto0gljpQUzsKQsE9vs+E9KjwBs9bwnZK58ZtqaiL0ZKLQId9Kt/JDyltE2n8lMehjg1AxkQX/k
IZHETEvAPb34LDRg0flrQPX3cwUDkk2jLr+oR5DTZ3B4HW3pvf42iHVa9Rl6e4XMQIzksqTKrIp0
bjdVkEIWkDgfd76a590H21PUoZ7HHgczEfT90hjbWKnFZVQnNpyVPEB2jJu8h6EpUgSDGwa/ktYw
Wd5N/cqq0ScEx6CV5zfuNpTfdEZeUb/1ZNrV722I6bJm094MXRxYDKpCZpsT5McjGch2DSfmyJb5
s3cw3Eyenn4V6+pahhKwti7UdrpczrjGMnNDPy4S+xfNhfg8VHHwvN0s52y3xPEywo/qWnkKKFzV
v62gPRmanXqDBNo5ysbmN6Slgb5jZGbP2PCDMaNKjDRKSl0L5gsuPrpXncYh3DzI2/rg46pb4mgP
J7sCwOzOnD8SQggeWM5GNYXtsg3YpX46jsAUbRqxUN0U1jFw4FaWg9lFlzDtD3x1Ioak6N6Vm7Iw
aFiF7AU2wQKi3gLKq51p0IqdsOoce9FOY3ibA3fRzugBG/icKDyOUxhc52Rsen7P+B1iqKp7p+g+
kc2GLT36vCmRFAw0Ko9SMFODK3qLaLG7+/4Wguqzmg0jgYGvM22c5yuzw71aAxUGfl8JQYR4mMPc
LaHoCC7wS923ew27olHBURj+zBj14yUGXrqtc2mJAZ086M+uaz7QXLhOJCrPwGG0SXOr0+YWuX5a
/0vMs3nZvsD/8tXqC/sGYVcf3IDpSvx49uH76fW/dOajkXfpSoGhW8uVGhkuDZkGzgclsRAuuLQi
RM3xDHNl0iMjdDRugYkg873R8UuLL2NbVhrXanYMdmma+bsG48hWv2bcxRdV+E0P0NovrODyaY7J
q52Lft9Fp/gCcW5TIJz07OhTtIu1VqqyFgvCJ7QOVsJqrhmI3QHpisDYIP4htqO0JenBBMSsk9Lf
Mbz6KunCir9MVgzXs5wkhmbIGe4HCdbo7SYVnEKlTZYWJb7eOHLBT3UNO3af+tx3M9X23yzima19
KOV7ac89kY6QLsxPqZJ/RzpsnilHUahRgNWoZqaXwKM+bs+ObfC048Q4ryzQ6HOoysKouB6XYHdz
6W3LbFCknmaWYJPoJ2A1x5u6VdszNAmh++asyEBvsW0luCjbhywqUGNKHCIMPQipzLSgscrR47ew
GrjFYMNlGK33ChRiI7ZPTXRHwKOKmlWEUrDQVF23p/GdAq8KzJBG9CWQyfro1hLwkcV1XdfLIUAp
9zfx2V2tFl13mgHkymvVFDIvjB4kxjsaQ1RYkCZfQkV6FWxhl9EEZrjAAilMdhfCRXVy8U7/+OFF
eKUudGY9rWyVYzw+JhG6V5fbaQwvPQKEDkwIzKwZtucCcp3vzwrDp0RQbV4hOPr4DszW6WUlkl5a
QFilYw4ZCqyMHNDVPEMMd0+GYcXAEdrd9ma+GvR9wBN7nooU3MgkGhJGWuH/9TcnnA/ZoYNSor0A
/9hQiia6NgM7Wrp9tNnTeJ1sMw8frrSnmnksvGtdA4oeeLMk4EZGkoMyaQfWZjuILzcMzeqGc+Np
wAy1OEmnrg2w00QBiw1Jr41v821GgZss6crBRo2pyWY1zKXfqWDOPmoUwxDz1hSs3ANM9Qd2/VjK
be5w/YGAHup05PB+abp5rno15yti02Ft8ypnF0lQkQMs+XkiVIuE2ylOHx1eMh2eb5iytdi1v0uX
N359eN33tMNL9elvwlAGc9aCx+uIqRyTzHe/4fFk/v4/Wckgh9m4aaaK4VwWSrpkwCPf4r5I6Yup
xZaxVzRvDGdDbKy1saInhCl4jT/pEHOgdKcXHDO9vTn4xPi0505DjU/hsEsYtiNl5+6gh1c10O8l
qOHFTSaVSVeE00s0ByW2U45PzBKfJqvbc5iUVnJShaMhwMXIR+rC/HHIvq7PDeuI2E7EYY+Nzisk
zfi6t/YpnKP89XSyFiGjZfM7oEqMJtNikX6E49pJA5KlzwPkXBFsVJld14pMuluQdyveSioLzF+P
3hLsRdpqFuWjpvAMbjKPk/YDBCSYLZZzPPVDwzYIORufJdhCwuPi04k0qx153WUa1njaCGrxA8BJ
eU+fm1eE/EOFiJkNaXsswYX9oBuyYlMmr2iwOXOMQKLtshwyZMz6Q2x9j2lbmNVkyDs4UCTQ5Mjo
vtD9NuZGE84yQLYwNMQZsjxgVF1q+k2uE8ld7MBviG/Un/4OHE/KpZhe8zAeBExAfBd/gbf82sSl
D+kZcB2vYA67giITje7QcGELuSxyIA77qenlEXmBJ8cLwUCe1dReCT5RcbgL1HrRfH3wfJS1j7dQ
IchSDB/wi8RN6mzIQ2Kn0uwMBoWMKhBTO51+TALOviBM0isl2ndjOCoo0Ljs0lP0Fri9QV5HUlwZ
acAfB7mKfPGD8JhGsFBKVdpq0pERNJz33/7ZOFgrB1KFkNsdxAp9lNmMNtDcsolxRs6IqFj4Sk1l
XBJsUoAqucWT4QI3unNqlNmhNUO12dCoGKyekcRNLc8LQi4FSqrUzcI5DupnItSNZcjdN5ZOgiiF
76dcawLA6CvTZBQmLrSHTT1y7iZgsmkOxHKirL08BfeYX6PHFXNYWKzrL7fkL/3xxqRX8hHgdNx0
n6SxdROlQkcaeO9yJ+z7IfOPauQmRmDaoKpZQ/lkJue/ubnzvnpApwjIwyGQJL2EmDG8toDm+E0L
o2DM3tNhk4B+Rp4GeCL/KXSHa7S+ZMmwSA4/nGrX/v1gZuSJtawA+VxujyqnedXYChzvm70E2r8M
j5ZRa8fngybRS0DWPPUYBI7yA4BjqrHztjP1I2BQUCw0U6iyhKaybCl9eK9bm+SySxrjLHNCTVkz
avbdANnyL3D2h8i2i9ZlsAZvH0OGanODw/lNfpIND7Lp8BLxkPJ5JZ9hiy30qTRkV8mqYeWGC2/d
mVt8wag4c1tAYcCavn3OOjdCR2jPNrt8c/YPkaoBMa3AWPqFBIwHR9hug0Sb8t7GhYzbabMhHpoE
Iu5fVB/zyDtAjVhtZdYoKBdOILDjouZRq5NkJiXTf9XiTmGf1ik1sYlOt/AqYTCRDjhtdS0F8nwA
IHA32wWkWTfypgIap8+Wz5lkwAs5loSqEw/w8XiAmdf0912trsUflJYDVWz8Nn7Z7AWu2KcjaItv
iIMgUNAuHqSzpuJYOh5KeB49/sI+zY/C21m/WI5wtFDXtf69xgwuhBRf3KuixAHm4zgpK0dHNkkV
xdMvC43eNR5SrsZMUKOKKbAjDsI1RF7KCLcWC+sq5TsJPI7ZvOVHeFyLFLu6X71AK6WxIUPZqbkS
3AaaFAlPjy9tn49bFe6YJ8GwYm6UTkuhH4SnA6IsY0Vawoci9m6bRkE70ro3Ntr2pRjSbcxTcro9
42wj1DD6Ga9YsEqPqsg3RkzMPZ5JV3jEvCOU4iqPn4wh0Zx6wK3wqVFR2y4gVADMa35m5i5gpgel
9GeHW1VnnKDwYY5gPvmw+mmzeT1kWQaQh7d0hc/jhDVrKoHyw0Ign4IEYmL/zpGP4hopFK7vu3TG
x4BeAUSxoEVdFMQof42BZkj6qMtBpmpRmBo42uOKE4dS3N9cDbmP/Dwc8e6YTD+z/pShohk6y+ap
8qXyGmblCJXXG2He4rlet5uqrrOQ1pZmGv+IrV0dyyi+OMXx2Q5W2AuAdUv8Ezj/7crQTyyzfuGv
KRKd/LdzPyqAstavLW7RqTOpU/43arkM6Ytrwy9N+yPHuQKpDfD0m2PDgpI8O2SWr0+EaILqd1NM
KBhBjhmkKMPWmq3Nu07t3sKQZZtvNSlKJ1HHmtNW6X0Gf/DRaxgYMf5/8tOqEj5Q7blqWHwvpNoS
n/M6/MpFT7wMz39Iub0B7GdatlE8fYnUGkOD3yBmgS6EzvPNEoLW5PGDfkcWC/I2FaQ/wjYE9r2I
hZtKv0Utua156HpAy3fQmAP2cFMpNOLtDWUEQLTu7Uh66bSM965iLK81ELtgC20urENGMKC5wZoa
jLGwa6UUvSoerh8NRCWEEXwW1UMOwVHuOCSHl8ze/s2w8GiRZ2KK5+0F0zrJVT//cEZb1wnAs3h9
bkPTsWUxTsG5MaybcW5oj5h7Fn3NCNrOXqEO3X71I4PUgN2bz+zRaN50KHbdiZYONbfhSpaoBtqS
h3etjTYsDC9bIlpMB9rxR5Ak5GTbs4KKOUhFEHmki6Y1pPPZSl+GFpS7QxxfYqlV7HH0ROKQnfXV
TDSzQrOhdYXYLFwG4f+Sr9O3JRmb3HRpUH7lP6gDMnsE25uT1r9S9qdaZKyZNKbPtRjnhxlu7vtz
vRzZfFIXugVv81Mp8dg0osbNT/qbGrxNddGAR+ZfLHq94MxRnNw8wjZqzCkE9CywWIOcjXkwkaIu
u1auTwQG426DcF1+CFELTerFjian90rM+BnO/msaCloWDJCj7sUeChfCj0/s8mn2vae4wRWvt3p+
Xk52F++5mAeTMV2vTBVn7tq1xi8PTyj2HcOp4vVTt9hOxgCjuumlO9cxtuL/boObFDHKirVPD3N/
QMt87eiGFgs/o2tq+esEW8cbHCRqiHQhMeZFv7rAK6J1y6f8H2+A8/O3e6ZWJUvZO9Qe+O7xmlLF
1ecvA81XFsNZ6wnUScKC3CEixnXWw7jYDzaR0AsYpz6t83n5OK5aMk1AaDf1cw39V1Ajit6DhcnT
Rb/EQZYehyUP3MLmcfT89VPLGEwg76rQCLBr2Zh5nfcjED4xUsDiLvXYmg6hIlCmu/ydkeibvsMX
wp+op304/BlNRf7buXW6wpKq8w8HK1mZnHOAka5O1xHCnuZFPMLKEUQocxudEFXpJPv2ktPIzSXW
dP5TGypngr+sYdBPfBq0P0G9+ACRkyO/w0NfNb5yE5UsDZVRTCj/bbqxuohIJFt/0D2Z1msSGDBA
lhb0It6O5tqJ1nIGOWbI82EUI2i9eIho5GRhM+CaQ68iUEzZ/+WhJyqi3L1TZmSECYz+bj3b239q
5YoxsDk5XybO1rQr3IPpZnOZzo8S6kMiwApgQq3Za9/1pSlS8Y7dVnG5RF6L9fZuWpqEZPtFu4T+
mq+0u7sWDa8kLe4AaspbxrzOm4pHoHmzIw4qOZvy7LuFVv1j4jhWMXYTjTNTP5dVTEflehxY7bHe
u+psQtnUMxOEP30Gk+Ww+ErfB1IzU/XiGztlT36BO80wexC4Y529ryCSM32OlmnbfXgQE7P5zdhl
o9KUBhbpwiGcT4AudJeuHRhLNv3YXN4F3tv0ERBwtcQx2M6Kgs7sUZ3w5PgZTh+6iKxJDJ5XfSco
CyM3bEx0JkraBjQxlxnUa3RCBLDEfuA7+hLsfQlIIe2furEbtBR0La+m8mgThJcMzz1DD7m6eDVW
WLoypa0q/lNtW50c9yIWWKgH+XoqwKNz0t/2i4qNMr2sdV+oHXS4i/NZ+tqOx52rzOi9XzQ3blY8
kRT5Wiy/w1+kH+ffVSYfQ3dHfSYJ7BMnVxpxwVRmnOVB7P0dwuq1nmn2b4oObCAS1FK/cQdoInlp
yVq3KFIHOkiCD1iEJ+0AiaTiFrrHlOYRtQVhnzs9sJJiKrpA5Jw3070eyBBR4UuwFzHbkVJhg1tZ
+mjIXwV57HEluPuulkd7GgmzyKPe2btlwRKl5rIr6CQoGFwBClW4Vo49pmWHEO4SAi/EvJPqYgsX
Ls9ze5e+CoY+zbRgwPhIzBU12Xhar5SPtFZmFDXiJUeVzQ20yduSfTyesqAVjYO/rkJfzi+rRArZ
ff5TBjZG/SN/rQ3mCFHwzOXRpAm/VBfibuNsCTA90GITX4O5cER+ulC/NiTWCh1oicIpuZgPVj0O
KokrfE37Qw5+Ff/DgXip1iFMJ7lWcZK/I93xa44qjA3uy0X9qEVhY7vaK/f8jeAhF5Wm/WJKoD6I
CLdPTMA1a7BUqhJtlOahkCEoHXlVc+8Ex3Z/eJqk++3FxvVDVj++wplNYpHiNZUx9BYUKZcPMbw3
8BtpbE5KX/sMdpqv+C5NiQs7PQa0uUAH+b87WOtdlbSAt+g/u9ph2TeXZjYcjZfJ1WM75PjT/cHB
m8bKWrTNoEDimyTG/2n//c1lXjshvXKmXVIU7WKXFIMF3KbIt8FClflKhXF/lXBmrSaFKUMkcVlX
6YoqgwuiuKFbKcjTlSQ+Z39OX3xSxHYSHO/geTOmYzX7UOZKRueqQdmA6uv3wjQnAuWd1tLic0ID
DpB9S7ehdTf5C40d+rUp2z0TDX6yEv+b6B+qFxIhGTwyo+1W5jxbQPzlCvhFxuvV2xUjZaFSzYgm
qnCN4lhkQaXAliI9sXmHSeqiuNIfZsBAGAj6AMmilnpSgxOugKcp49wqe6JXDj9cvidqcNDW6LbK
dtQBzFuBqXvOe1zad52oBUTdfXBO43MCr/7yUKaKfwzheyjs4TYIkippq8gv+SU1i1yWxApMkwNH
Mf91XWdoUfGCJUmRZnvj6+cvV7K6FD8oDZhtHGRhnzoQJb0kFIWV5C4EhJgF0YWzmpv4OTJ0AM45
rpt7fnPAoCQmKOglSMB3rMQjFDNCkqAfU20M9t9yIJESC1DFF9UzaGUKeFmkJr1MYPJR+L7DPpSD
76WCyYKpVqR+hjIbdRJ0SR+47pcfJVISBX5uIpKznWNA0erUp7HVv2o1hmSgNiOuKUC9C5IKcbZ/
6qymazo+muXODCLrduqHMs4GQIF6aCFwpIuY6Ay8zw+QkK4EbXx7LM80cyKzyJeS+xyUVvz91p9P
E7PTfQDMfLY1ATKbQRGbXrM2PEwovv5HOhwXI9qCDagn4y8+7hDhIUqpcvD/XJoM7O074RXF2+z7
NHYz1sbrhKxwpoiIGdV4+R9SHFkWPo6g2sCCsfwXCcS06axuW1iVVQl0bK1VBOB7jwnAHODMnPhK
r5yrrG//mjGdPE0ID0u1EzI8ULHBWpmSjpQbVzmquJ3nuPMMNPUojp+8MawG/b1x2YvaER4lNMWA
4Px4dbalh5dBGmJzs1Uz4KgEauLPd4TnkhXvOcy5sivduGE5ptk636bL9lHcQK/rfmVbW0dnnW/D
QwWAJua6fRzyjEVtcencmHCeKL7LoeTJAm2MODN/KhfMUG6CTMYU6/01h1g828dbXuN2gDofBWXh
E1riBWCsEPvRonvtfTFypuqRuas0p81p1M9uEv1UFOkR2l6iEa7U5lr+UxIs28FxPZqCPyvy7p1m
MYWRtOTdEApNuDLe2a5C5IDN/dB0LR84oYn/IzsmPEuOYTQuPH0P7Hek637kmCYhGnFw7xEGOxWP
XxmNX70w/Z50eTgzQ5zlBZ7vh5DGKSwVoW3uFfyzdFqFwuEMdv11xQxLjDeG8p6BRq3dxh9ryMub
nH9rDsyg93d/k6P+6wbjQxhH/fFxy4pRuUuQsiPJQWmd4QzbHI6+KMXWff2erTyuLaAyMwPTq8er
WLvAKZbNCqNY3LieZMDm3r4B+3IgIBB+wW6yK5htIXyRK4QGLjYQ2SEsjMkhZRUoldBQINNrm9C6
CsOyJQgnJ6Lh+92nNFoQ+Mt9qCcCEoYqZ2O5Lz28LvH9stZ0TRrq2qOxGoU1aH2kLp0VAjqE+WtM
OqwTkkAOnRYyD9jw9Hiv8sbCKYhL+AhCVSeEDQpbqdttye5f/NF1YjEXMfFBLOPqasjQyAdTgPu4
vx44P6bjwEhgNodN0dEcgszCT1h7ckIk0vb2FYmdBd+BqDVXJiZkKUh0E53x0ISIrGu4i+Y3KYzi
rD4BsL8d1ZjBZ3ruC6sAxUtZRLkgUHmih2gvmc9YfGSjsqI7qQebwwqaf1ph6ZGuapHJUOo1t+N8
dt6ve6MkIvaFcdW639r4btYe1d1VbKmT25BuDOsLPD9e5vIsQ1APtgKwWHGoZ7+mfwH+KCzAAlMf
+DH6J8oJjjwqhSnAkaTzZrm/2r0MRyWW16FfuMFmNHr/zJrG/Cvg8SvdIT1WrXi4j1F1rfGOMd2z
v2Hm6iMjLvsHgZX1ieGiTQ+AvVxOAsy+QqaMlUQgx1b9SiE3bmOuJ2YR2UvL19LjhY6RFAQ6p0uI
eR+ZkOaaBpdVzKM84CEAWBwDnZqL/R7b5aDE00q1Y4zkqbPDKaCx+z8Q6Psoq1qL+FzmcHqCeTCi
whQLmBK92mLxNJ31jX2wfYD34+PYoTsoNty1AmGVFJDJfX5H9ofaT4BB4Cf7G+y8RQrWAGlvbwVO
lAtywQi5L8MKnGBsUSsuKeIrDAX39S3q5WNFSH93QwjHycgqx2PhK9GpnmoqlxhTNG3jVU1LldOo
o8UrNYsHcIdf0b+ZruQvjhgf3qC7zL/4NVISjeus80xkeODY4tBKntiTCwKP89BL5fOci695Rcuf
MyNuS3VvvKMyZchgaA6bjjKfgf3ReYmd9nhyqOIGEV1WfH3NfdZy38nN7HYbkioqQKDqRCDWYGvZ
tV2PNacyIsY/vf78j9dsCmSaJN+agBb0j6vRABFT0PxeIP6Ox89j2sX9L6H+ucQ7cyMEY5OhYOeR
dDJchzlHYWJJ7juL8SALo76Q8ysQYTYS0i6XmVcOnQc+tMmgk2eXd7SZomHoxgDd0OWiJkR0xbsZ
T55O+frOfWXr0U1U9hjlznnZT6nYCcsV/DhCKweJ52pw1/VD+AsZ6UjbotqkfdGCHfAKmVTuTMux
ZwUMpbdetC8K0zPWm2/buCe+WH7CLsXb9tP7Ym8ghBw+27Oe4JIbzlX1yj707NSn/e1ouXEeDMRD
9v0/oGVx10XOSCmjd6n1ZYhmnEVTlkc+dgxS2tNcgNwC1t6XsxAWN5Sh+rUWFXQsb1NJUS1SPgXV
LEgr9D3lyliDUIo1uuGh45x65hId8KeG9INav8KcJ0W9TO9JsZoJya9Ox7WwViUAl2k7Ija2r++o
jWVu7Hksi7312EEt4yaHucFJmARx4c3Bxwci0RaUG+v36XVa845vECoSSvyAhkhaBIKCXFG54mhk
RduNbKtnV+2Ee4wKE9Z+EdR/+eHzRvVpAdbG0yx/p9l1TemWaGb/O9phV4WzDOYbIUcg+RJsUDqY
3zD5C36hgg87KnQEJWG9UcJYKVmSu/agJnw9v4PkoB2Zuz0mXsO/Y6be+u2wVwLPMMbCs93ayjS4
1tGyQdkwCBbhf2cAZEnu5d5CDgkahmkRSwyEUyl1fRaTmWlnrDhcHMjgPR0Wfpf1ZDdKFR0tXO3O
N3syex2hidqfgtk1jvmK16h6/+BpZt6b8t3V6amx7FNUtxgIRV8ttmxn+s4YIe7RfsOFgy4HSAEM
hL/M8tVxyft9pDQzt6SpOISV1q3SwHSv6kxWupiFk0SH5bd34RDbqsLX9hntJnQjGxRxyjwe53Tz
3Mp0kE7t4xhi7IamoUdv++41pACTrkapumYOUxte6I31tF+wZ/D9TbfbtNkKuKhvszdjZcxLODWe
wnSnTIkFuErM9+qOXtecPEYRBWMC4gf2PuPJnRJVSSkBwgYjAIjyT4F5zMGX/og7xbprAzYSekJ/
+mWC0UI1gL1IMsXZO14VcvJky3UfUFGnGcZLfi7EkYpYxEB37Suyjo4NbzqfgfdZ38yu3lmIlwL+
/d2bP/l/hD3GG5IsNNddvFVOE3U1BVpiuGm4LYJn1yJtIsts1ZNmKPXjC9lvK3tXQ/EuimtIpuB4
1MqtOui9UQVHjd+vWZBXNNM3ROJ7vbbDuz/W+uZvXYyIbI22/Y1YfCCWwDXLQEaTVqwfdR21OwIj
b9YSLdn93/XVf7mBIo8d+gzXH0n50YFfnGinSQaZIFnO747XOaxtc9IqVTpFr+ikSxZolWHZ0jDa
EZYNw7KMxgegXVL4dUjElpvIcgnOSeqIZmje7EmJTPSTkxGpKo44GaPc6b79AoGMWKm8YI1IkWQQ
+92F7BROTiyc1M0jc5vigHvCKpzCpPzWXru83fVIxu0f7j2VMlJUGxYRjBzxlS1Dqht/YWBH8smT
7UA8x4ZI0iW4FWcf9gtHUp0/LJX8F32MLOxNaiwUPOvLMrJ0/dRI+NGRC7cPwAJLfUzfxS+mTxUx
a6z5Aoxej6K3tnQSxs9v/iPC0J5uWz/lgNr11zYdN6tIxsKaqChQt1F7If1u8rj+YFJFvj/W0rTT
/ha87f+owmGAsBcZpCnb5mLvr4vhz3Z833T6VBxufwu2sdHfOXoFOhZH7BmxlrVGTR+Z+kwSs2Wn
YEINy+/LMVQqSntlUhr7cTdH3k4M3YdBWGxUV9LWig3g70G/8yJ8iIZDPahYmL3NMq1Hz4sMusBE
RyF5Wt67L0FC5q+40YasrQ9nVK9V6PkqazV79pXGg8Y01I10Wa12dWP4jDK6ylFWIOYa8qt423HS
dIhmgV9fMuI0ueX766yx/F3RCqCuTPKyPKAS/AMUVH1h0eShNrSyTPpF+mTfMhr9VS4gFu55ekMo
aoE21JZ1EFdk6rRIw0HfxRwAmZ2t7aYKThYfsPpxlsfEFs5cC4pZTT+1QEtVLCHA+/qYAluR8YDJ
Wqb6dRnymQkBhNVn2VTIdwxt4dF7lZJxoq1F0i3hh2rGp+CmjAtwZvRW0KJjvOOsRyhcO25zIKVX
r+8rURMlVMbwfCOf4C/EtLiaG12si3CAu4kndenmVRFIsFX/vvKPR3XrCnkUCgG6uG4SIeWrtrJy
zzzEH4Bp8RfMd59AgHLNZ5qC5RTYyA/I22I6Z87NqnDW5I4qd2ZWMQKJrEZmPaFMprqUypBDgry2
Nh9NW2EczZJLufYC47FYDH6qDU/5UHyLLDcMQuZ76iL43Hgpxsy2LpkiMIWVvVYLO/tZp40D1Wpg
xX+dc5gqZKAM4TJGv/jDCHLcmevGTvdkVysPhiF9+2YFNTH6vCs0D+v2qZEiJI4X8uHNO9x0ldzB
1el3TUQUM75DRf7pRXq6m4ESEsirdSKfU8IWzExktcRnVIgk3YwYw+/bnsbyzSfdWYOzWY2Kg06C
stkBMR07TYyr1y2yhGkpxixy3u7mtXLeb4Okx+s4Exnxb//zHm8O+ezi4eFzfJHf97KAQVQZXPhV
LW/3mL0gPhloalFo6R+3LuTTtntbGkh9seLSAdF1AnUPgkalCM05jsdapooRA2x6If1YjzExyRZU
mdtDto+rUpl1YKQ7Cj3y99cVoBdTfH0X12kQJZAcs3n6T1LHgPpCzDml2x/oUCnXHWRr1YQqOKX5
CGkDtJA/6BI7u2NjdcEujOrb14upO4RelrN67VvAQDDL98z43bc+9vuny7+u6hg7zTrh7utyLIVe
VoOeEcQ1DxmJ9lAMdC1zRvDVo3DKKZYJmddAydN4i1OEEz4CaGGY9+68M+d/AzsX91cXBbc+XkPq
3YBRQPzrBE31NYxS1YAMqPPfiElgSmPzB8lKQTowWZ10ClE49fgFFYWKuh9wa5A8ZQsJASeUX1cc
07seETPaCu0u1+fnG8sRbXsvsYfk2RtvG+g5mZlshYZ0BOZoJhNS1xqGDTItIGOdm+oiNw1PZPra
fZBkpZL/y4Zq8QkaW5xs9RIjRz5yTCdH0F9pPIq7tdku+jNk7whxo/+o7t9bc2nc2bKBFr6o52ds
S1lEnx5kPwhxDevnefFba9ofs+NQz/QXY7I8+yU+hRl4F/nlrM30tFYhYTEigCMXIuawZsbqeYmi
M6lBqNk1Q3k1jfz2uGSZ/aNI39kkkNjmTGvs1jUuG6it3qodb01vv9Ux3xhKXlwahjyvibtIAm4K
L0wVQL0k0Q+i73YHDZSgcFCl53TUOklvOh+f6bqeePwsycnuU7dUcFGOC7/Lm81sHYxZ52BwGWG2
UGWM1jXfZoyOt5YnoDShyxjSlm7mHYA+tgSbxcCCYD6oItwxEvFTP7jbMtg329v5FDbJVWe8EYBO
6l8+pRsukCA7WP6LjU8lTFiQA2HubwlhXlptmy1oUwMGgRUMmQlzDpjNt9o4Soe8aSlNT+TnOL0e
LdkC5SQFrt1aEI0AmK7jrFOcG17xGPj63bkADgL5M1sVubymY+ItGHI+H+VJpaTh9/YoCvty85Ju
T/0e/b9tyBCjKNV6yRc6QNwBeHiooSyi7qCH5jby3uTGbnbr89iIgEd+FoMaTVKM10rQXbSdlHEu
xZgRz3un/oT9PQvRirxnhlpYw1wvRXAFv0Tas3C5MVIpz6gLsYc/7LA0lmHFukB3mWnfED9k44NP
LZASfgU2XCDaZguuRT0MvmrB2wUf2uyG2MIjgMlmYpvwpVZ/12eOVqItZ7tA7FmOJLDpzfVL6v12
Vu3VmPlN6vIlL9TfeI240n/yuv2quhBsR+LGa+uZPwTPSDjbq6/RLL92wA6grKdd4IWtSnCJ/L1q
aWA5fCBOQVl0fSCWYy+2aQzB19sNS6UazPhNwp9+CVU7htMZMSxP/gsFq7k2o0PX8rGefwRU1xRE
Tt/y5Pb9UK99fmLwrHXRmWJUWJTT0uVaITqQrx0dHb0lG9J0U4SnrLfr5tpRJ7xrOzRqSLKqrEQ3
QgV8JcEpeSQVbx7vbm/UjSeDCkkyz6Ay0jLZRNfXJKWiP8Q8ze8/XP7bnmiQMbURYD1pSGerdL/t
QD1xvdaDB4vRH4CPz8OWHyE+kBr2EJAEURvi8gWvC7bgQB0NqetQvS0rQmZwjRMzF/K/N98aDnkm
dw1qsjAUTFHd/2CY3VKJM4RM9/GjCQ7G6PtQImX7j9FQxIvkK01Xrlu4nBUwOaSlAqMzW84CAYlH
mojDGgLeC/fD4vCzm9a9PrvgJe9+uNmrWPKO81079mYVJevMZYASE5TyCPaW2oQScPHJwbJ5pYuz
jgfUl9F9Yt7Wc1q+MOuPbytBB+wKWqBRtPj3VxJTR8X7hvySPt+mnb0k1Le9QyJ4p4/apMHcqysv
NpjPgkwyC2+DjPIcr7j+1nAV7ZoJTdpTDONApUIiom4LXrv5B0wsr6woQKgXJiwSMacKY3iZ+teM
Qd/dBiymHX9qZuaJ+dNpEUeuG7EPGENCZ3+QVSQgyGCjVWunkE8IX7XqM1hJKghnHRGhRIscGKvl
3D3NuPTbFRlgfoFK/fv4ETs2ACxW8xLN5czmxSC6jatdHU0+wTqF2yvIH4nvi/UW7BVJqlcQA61T
4IvUUz56oX8Xpur4EPJS5QI376nNRHzp5YjzYjpqPPPF07L7aSJTEkk0cFA6gHhPZ2cJikzozfPT
tbR1EAeaMqAQEYw+CfMVCwRFu/60/sz5aLO7yd4EbDigAy1lKOh6KIBNDNXPxvhGB2kbozxdTLA/
FUrjRdc+itXXqYlqTTmqRSVFCyuLl4frNeBFjR2o2ADyAz7C1wRUuTSIWY+P894qob6KXsvtn7kn
WITvwPCDIX2QfaJhFz4+TLhl3EWO5Ch2Jx0v8pqcGJIjOwlSKTfO46TSEo7iyzqgqApn1Wub33jY
lGNlRjXLODu4reXyfzqJkqoThh3AF1zjDNJU/KXR/xyvF9DTnXLaLz+xm/ppz+IzccqNEj03Cvh4
hiwWpwHSPwItod0UFmaT+ZJvu+SEPBYPoQK4vl7oj3PauorcNSF93KPHXaseZEJY4A5Xc88N0juF
TPpfGHAXTRI3TA6gcgL3RmEaP41P4+jS/mrsVXbZburkRHG6xzFe8g/1z+iCKM2q+roRxWSjL7B4
iQxcBGMMaDxLwzc1bdzoQ/UHV7vCMAgBszrEhM3UqmYaZ87ecpuqhHK+nPeChnys+hSXK17nCTFA
SFw/P1YQwZVNm36MAsK4sShzd+Np/tiIroMrVjRl7GQMsru+2ubVxwZwkKoKBimm4dEZx7NHF5d4
XWv6W4tvEmSixXklVARjuxZN7KHrmktnV+K/y//bfV+7sCGkTILmLHQ6OfmNwNp3vevbTPboiVi7
A6uynMmMBVLxVWsoycgxTGvYZW53jzcOatTD6viDwLqfWJmNDNcW5YYO5hMc1T/LNjhpu75nLBJ+
mQJRBakLYF8SadGiCLwof8Vam1+GgFw5g2zWDEtHaxJSb8YM69qSo35TGxYGYwGLS4o2h3O9gCM5
+sNGr0OnEWv5oRQNPv5YnyHYVEto3oHp0DQ80cIJgdfDZ1tlR/p/wuAP8tOZgJr4dNW39k+r4TjT
XxEN757kzsltWzXCSJy2Cx6yyTGwiV42UKdiVr53HSnuGyDjBypgcT5InnJLBj7375Cok6sYq6py
/YeIz0lXaT0knh1ooT2P7Gg7QQd8S2BWDZ2BZMajlC3IjFGuxxDHBYZXp6JLBRvWyMx4g3mUkQeB
oHtpo5PIsBjPoW87ObvAvgcnd1lvMpAAD2i6hJLzjP9UdJPUfg5vcu6VK/gk83oElB78jkCdL8qp
2ezDr//dw/rmDUlLkuheccIwVJWYF1iyFSe8s5DF2uBUE/7hwSB8vP4YhvKUfEZkeRsaxPDkOyZx
J/QsICRGWLLnVAN3Lc2gstaEqjk3jeHyGcnHx0b8grFb+w6Z06+QdRgEDuZXNM6VT18F3GchiKFQ
Pdy16yvnu+SjQ/voWnNqeGyob8rmXAAViJeEtI/9oBVbQI1liSFZDokkCcRz8hublw1+BqIqNE6S
o9hOHnUh+kLqUFE8EqlNKzC7vRKZj9l/ydNHlHrquggvABfY1Y5YyxAEgZZB4EBfGEVXwdJ9hQNf
aZCTd1UhUs6qVlT2OhO1KJtiStrgG4A6BgYIpjIpwPq9MptlL/ntwDg3JEMcSSofo0/bn9124FQm
BAyWeiEf0m80Z6szezOvNExr9xmjWijz6qxQhUDvJFsQbbFd0Pt12rwI9SmaPmYf4di9IIbxi0bZ
iUVqMEh8t1cfZ9jxEWcaTcGvHuu9/K7MatanZh72IGAf4HLyYpoSpnY363RAGAW6w9Ep4utiXcZp
M3VA4o4pnMpsUR4i22xPt1HOyaL/46x9EKZYCQUErH5FrAZ4FKn/RfR7Qlm5WflfgKgWwkEAsd73
aagJSDIEQl+x6P/P8iE6PSOKRS7MAU/2gVv2R74wivOHja1kN+0lA/OCtgyzyEmMmI/bYDZgvHCJ
pF13fWeOskLplABhkrNVyknBDVal1IjfcqP4FuMO5qfMBT36K7D86sKX7KwWWILJ49Xjroi49tbq
txQuwecWSqY51f7KmiqEFofNLDY90j7F+4GmYwxKjEQOrcG5mISxjEAe8ZHlr78ivrRMnpiqGi+H
+12wPXux1aESMPGXmZGKub30+G6C2i6ZotavMZgpXLNThXoT+5lXH9hK2ObiPXyIJ/sk9I6rwC/i
/1rdYpuUBADoOwsmnc4OZ4V5HzuypWT1yxiyoLTXl8hKEJ8czIXAJrJkGcA/P8ClbHQjfSgNq7q2
AOu1ywpAEFqGCPOP6fdFNm+EcGO5Uw1+zS2U74pkX2LEPb6gewHNRGqQzYeQ/0brlk1SQrQ5ZNO2
lCCRGsGFK5Ae70E5HmIS8ljEBkQpxezBdecITzdNH8tTqM9QDOV2QqUFcWmRNnp3NLi4GYOCna7L
hzOGYzjAaeJD1bSkL5Wh4Y+bS5KSXYnEVo60D8m9UdYJCKCt/VIZ2Qnl/sKP4sCphrCFqKOmCknR
zbEpfvPk0IEAkoIRGD849cW5LragNyeo/I/vYC3GD2248UfzWwaVB86MmHE4/eURZ5HTEuiZCceY
MTpkMJkWSf5dKJ7C3PwWh+z5vlzGX/m8zDMuDXNF27P/lIiay+/ufDJrN4Y7JVtoITLPXFfjof4G
UA0jYCQIyJWrqNTnZfK6Ygx0xNlJNJ9bMlZp/L0mpLuINmveBGA4k1HOl7jhbmBHnxPgD8rh80W1
cDQpWumaepaeAw/e87dNDzDfZHDIRFeFgZ/V0gg4v+AqodD+S3GX3RtDiszD8WntTnupAxJLQoIt
zzzFANIPqsEwP3VnDOtPnqZV/nDem76OQi/GlBnWJ7jL6BL2q86J/hpTT8RBp5OzCdxiH2G3BRPz
FiDlKMQBnpeXbvjNNX4h/1CFaX1PYKJ2CxiCXV8E3xv1BHI7rsZwzF5oLs56ZemS1kOhaqhxv8N1
KIFUmMqXLmPm3NELvI8TPgj5/am4S8hT7dQzUQ3ZycwM/+/M874COaPPUgkMmGV1DJ6sqQe6UC3t
m5boGLNhCzvF9pwS48e3wU7rt74pSSDwmGpKDlFHusYkIdjqLjNkXcuC9JUfZTZNWK9woVMRT244
MRBFi+GPtBZD3BQam6A/cGk1eObFrzHVmGXIohKpuk3SgOuhgyQ3X8bpbJPBHeGKy1+VprVQ4yqE
EltjsRztzPE3za3Yz7SSya2oJelDuTDBdt5T8vBNdN5nAEC2k+6U/LY2Bvr9yRTWNAIvYaCHpdpF
dlDK1/g/C91FValX7h1Xp1/mbGgqNVV6/KZa/jO6ypVBgkonbE41tOK0AQzqaOQvIiiR1dgvv5Ge
5uADXL5uEfjHb2hoCUZqNVgnpeI8zgngZgBBczNCgm8zXcBpVAfW8tr956B04ZFN+o7mWbqb6PAa
WJTwfwhZlRg5+rrc7aQN+6kdhwShaoJQoCH3Y2DBAreSD5h4oWN+dRnYgGt0Ytgztiva3PylLXps
CmihaVpUlqIHG4WGMhmGFegRR8f9YVhAcuoxKFu2NTF7soqc2Gg3sG4Ds7rJHO9+W12gai/TBmXX
csiis2NCj9wp9GwT7Z2O9lEnLqoi4qykd6cT0UP+RcrD/N4/NAfL+4tNkBVDLjInUkAcZW8MD51u
orLGPl02dAXjeghLkOuW5ehDumLpLxqpLDOZsFWqIuxINqvNHwc+yi5bvPqIWHw076Vc03+6rnfb
FaO62HCIIO2wQQpjZcHQULNGAFT/tNRJ0WJr4b2dulYiPPYPPmWN0AIxejM99hm7yv8TxkqpOECW
AqHuMU7kVtQAKQvtjMRlEAlJtUDju0EcdGVDHHsDWZV/c3+EqH6Cep6iO41YSZk2MwWiuF7QkzS7
ZR1ocds6ktWNKMvGTMuQ33Lp1vx4ehSzH7hFJdhLP5nU9FQNdDg7RlQOiTLNSpqwsTvsovDZBJxd
BY7PSaoMTryVh/1tHLWsKosj/KZ/nyJlDUcNKztKc5PABCUIl7V5xHtkDA274xgTQ2wu7GhRUSr+
Fr4sZQMkS+bXNJnklJlt9adXUNvoxTft4vjCqfnzNvB478OZkFF1hgbYePVM4zqUBdfceplW3rJR
1cIgjIKQH7pHbo3ZXCb3iN5o9/7cDXp3oAyQfXVqc6AG2qmr8qFkIhfFGIy78GljoBBeTmX+vkU7
Ilo75tbo++uA8twjR1y9JIVcr47T2UTx09jn1Av7X3idNiN0xPIJYmOVUu7g7No6QTl85IYQJ9VG
icYPtasc5t29PAGfYVpHnMnLBJoG5NxPMje2wo6DBc0nh08Kcgh28DjrOn3PLFLsZl+gsnGkGVlq
knvpJgLd4dLqKDjFZwZsteuJeCme1sM3mncTLG+bIKNjUzG4ql+fjN+hcfKyDU1aRXilb4JymP89
unQl7AVtnKxVFygswf0ybRNCM8VeN9rCvBuD+2nRjhGGrxkjekttx6kiLUUI3lbe80NhZDrduPb2
JFB0QNRX1q8SsZxhqcyAR1uv4rUsYjlqrZt4oyPrZpw53N/oIkIAtqTIMWFzKFy67X+VeDfhiya8
CMBjgcjnTsbBXj2/Ju5UaDcpqnKkeEfWYCjLzSHNih9pJ0e3jhwmqB8qi5jdO7Njza97Us9I/1qU
TcVnUqfnjzu+kNxJ7pb9kPbZlx8FCQ+sygS7R3z2kpzlmoVAF/P7TtZEwLQbLsoJBwKD+kKeNf/6
vL/pd9uI6da/2NOsuLnMa3bcanhECAwMEGhzSGlWF0gpgD67mpJN4BC0MwrvAFByjtvDlbpK0P6e
JMcXQ3OXvovAfn4S3iJDQfnb78LLW7DUokWWuA5sYZTZpvOrMUOvwMk0rPV2qAac7OSdRAEDYjow
1nEwn5QXtfPF4XHbeEGCXBFiG1/QbUw2pv9BRmL3c1E9Qgrd+iNUTEpA9KoN0NoAlAf47du1YLT1
BmIcW1AOUdDE62hmqAK8g4fbKHS02Pt6hczVLXNlD2ANMxJWZd+x0sY7S4NqZ1cHNxppLXgU5n2z
2kyIsvnJkgo8M4BdvpEpXcMtRD/AkaynPSXhHiZB8CSUE7l6/aAHGMMAGtvXqrh1Ea8WrJlGpUbQ
i5hLaFOHlG/lbkoeynGVTSrvabi/w0DML3z7pkr5NUCoppL1u3/FDuE4R85ulsYQy/n4Q9Hd7qKW
2RLl4c5Gqh9Ak7ij7HZCB5IHc8OX18aN4E2hQxEpdNOpIS+TkS5R2sqPGEufXgoAEOtD5aMEycC3
wPCjdDD5apa2NlfVND93ixc4SfDh5E09SSWJJmIOtmuYCfGSmIWamY4ScK3IpDVxaIDs5p2naMhu
fOk29zugudVGqs60xQUW9qUO5BY/7hl1ngCaVMLaHEVhSfgQp7QbJpY+WBeHiigoBlBto4igajub
51b4MlHAyRcfnK83
`protect end_protected
