`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
fVAOf/4aRuOo8qbJQH7UoRlQiOnAjbVarObO3HkQW6Z2X4MU73JIB+Y0zQ8sg5LSTGExe8E5zEbt
8Um4lOIaRQ==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gJfTEzqb/sa5TETU3t5+9O4oiM6EquENis3Y1S3d0H8G78GjmpIufQebDT6zLZBUO3YOPfDOZpcz
6d9TgtLS0Q5MQeSh0/hF8AtmBJ1E+FxU0Rkjuk234Ctaf8FSoDc4Fz74AdyXAFnG9772oLL23oRe
mYIObSXzI08ti7g1OFU=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pjtjuKn3N8xKESUm3csrDZ64rLx5+dRzIwNsSDN/PpwKMb6G01EVdS7duiCt+b5J+O/RhwOSUuJO
CK/ix+StCIXb/LGv5u+kYDqQBCpkegyfMy2todIAj/E0P6t6fY4ZmqR3frq0AdJ4gaC7AxFBOf8v
NdHcCAXIq8SnegCYYPZlDuaaiP3LaqMO/F4+G8FS+SD46uNaVhl7cNKUeZmZ9t/YQ37kFJUfBCeU
XIjTVmCEjXl0avPds8Ul772f7VzRBrGNQDl4JduehAJtHEpkfej9pvvKoCKnfBcZReWUGyPQUHW6
6qGPzMVcgBSjgW26YvbtWuL+E9FdD4Pu4nq3JA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
n4n1xWrTjHv6gPz9522r+pNM+qOEI9rmIEKesaY4UP9lBYm0GOFEC9O3m0KVb9V/T+NZy1dNBsLB
R1J0YS32gxzDO6Sv5d1CYpjQJRtWux2OHLTJDc4XImXlAaRS1VnLgIzlovWRJCtVsCMESMI61Mw2
9OG1bKY0ieUNe771IBySWr5gVm2MzUkQiZuM2kF69etRz9bX6ke3EHIoWAT+J+B/qSuH0T3515s8
9ibLamrCcKyMdohTXIvWZSHu7cdtO3W4hdvLopcHZ3qm/Tl94UOH8QRbzy00hui+P9bALB4dpLog
9Yo5yre09Vl4Dr5lUZVZwkuTtUrh116CsR1DfA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
h54kW2YmiecZ77BnHdVTWtiySHRhKfdHEZ8AT5mFPBnMWeE4ATrlsYEyUkSJgsBp/Ryp2OuOtLsu
TmvWQaBwzr+Nk0bMQvo1ixQbs5NVK8xr/nFQr+hMEyq+meytgxhNb/Efn90gpqvz/CfQ78gCez7G
3AAAR0AbLGcHn0mEbhI3JRZHOitwY5u/aafrOlHqcSzThxa4VbsqEsemwTZV1SiRumoTtvGoquEk
eiLV2PkN7Dm89nQ325QYm8ZO5RErAjCoj5ddREby8RAbOY1vCfyCU8uLTNOPdWpsCDMUrF3hXyGZ
SsyVugrTSUzRGLTZh5b7xUFbUmQcxqqJJAJtwg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
C++ciYZRz+8yja27sV6DNrLlC1tZ+kZHi05eyrD48tDveC0IENR9qaLp5JG53Sp8Vf8wm2qEOwJ/
Cov6z8lkhnu3uGXc03xj+oHQtuEFnabbilyzeBOEregYolgPSKbR1qCHCG2IsBm0XohlxD3lw/r7
ahsJ+oj1GiaQruax/Vk=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IaALqMhvfCggMH+G6/MmLeU3Y+HWCFn5yem7KyNipfku40f4n4FPAGbkWmL0L8hyVUhZm8pQZnC2
rtcTwtFZOCam/iyOmCUCfUE/D4HUnNb1uA7q0zqBMCc3cbV78Arn+FCJvaSO7ylx46urNuiFfLQ9
TitTGcG1AlOOeKF2RheWfK+QP7Kj+pAbQcas/CcbJfh5OPBB6TZS0CwQStbQxMUnH5bjvL+wWyPZ
kKyqnarn6324BchqMpDxciQGuybA+WRYOv7wAw0y+Tte7tTh+5+hdlx6UsoL7kOHlWms8rxLLnIU
CZqUNUyORPsC+BchRfkmHkEZ/F+T0Y9avEUUJw==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bJFRR+6VFNUNvQQv3qY0yC1m3ZjbUq9Y9x0z4De7/9WMzaoWBmHihc2XRRrh4GljlaDuDgnl/Klw
S3CnQbtinjE0/o+Y1m4KCJUwLURuEIgiUtl+z/0YkYKnOaHQixCYKtwVrEu505445wbCHwFQ3aOG
vJyLZVQOZ5PdvGLYz+SFfbVaN7KaIBm6q4HfFC7uHvvIiB/5RcBMzUwhexBEgHmijGV2jxgqfYHK
2cMj2S09OKfWh66DxxqNAcjyNxpnmHO7jOcCA/Bfj+lhc3fmnEASd+CpW13so18tYa4E8gvLDeB5
S6LVwao1KR4Wa6lN5GeXhRT2Ru88VADwofRXjA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20128)
`protect data_block
Nuv6YW5RofoA3Hpi7yTcfergAZI+BWziZRxuJPfHpgQ3vZWxGgnO6tvFA8VF02hpq+K6xlzMscCc
89Uwoj1UwfNvS4i0ZdeAJBK53Ag478T/GDMZnBaRoOicA92yojt/2ytSu7POMpREdBrvPYK4IlWr
Eh9JMm6ohxluJKff7LqEcXfWTi1El5ccM0lfnrBSkxNXanNjuFUrhoCBD/PwApnqR2gGcgXHrRMx
IM68IZ+NQjY/7dLTuyzuBNEOe/Bg0/a7gEktX+C+ZyvADtYieTfYNJ9Ebk9guboBg0Wx5xhWy+Ul
bVHXg4XZKVzTwpeTVOTM8ih2SyY0g48pnJ2xQzE5H2frLER2NJSI4lhGEcd7RW5TolZwJmTpmNdG
j++fviWVJrhEECpbo1YknFVIKK/DoYueW0gv4GegdO8stcCdDjXPTkwmvbk3nlVHWR5LNZLIenmv
Js0VnHjhbQDC7v+ePKf0tiqBUCM0dITJ8QyF9bFov5ofMFHPbaRpONLz/T5E6/1m8R4PsCe+AMpJ
La05DFy1o9PSjW7i3IVIwv1s9Lyx9omC+f+N2q0j0Mt/OZe++OGBiGrz0scBL21rMnN+86zNrVb1
jB9yNx+1i7SHa9WI+3xeUzQKI9qjt7LI9wFz/61TILohD71Kv+Kcw4uV+zL51jyZGJHKo38teVFo
Rz9KPUiVa4NXy61C5KzDs/xUKHZKFgMLPMHhj0dH4tAVboDVHRbwRZrD7Nl/yGTix1UQJZJIG7lW
j218cjwSdEAoTpx42Omt1CzswOVHYMOOE09BjKEGemKfTUqD2orSMbl3Tx/dcnoF5wxkcinFL1o1
X4ZCJrhDXHxudN6iaOdeHySVcewLpszoxoKvNgcdVrsOKf0viPnhmi90XOWDzLnCRydE5zYMH1Jr
AhspClXQFfj4IQs2hM9XYO4d/6DTBsSKDvMQN96cP64jcJH6atqo4tCPmwzKmPMY1E6kmzdFWvm4
6mkxnuVl9s2Ro/mBZcerDvbvr9tG26eOlJCD//UZAO2zNdt4Cha2GgdY2ZsrgEj4hjEMY6FyPjrl
I4EylPmu2viOsEyTb8GCapOaYeWWbvIXxjpcwXbAzSe6S8650SYYNbZ2GEc03I7dtLRKOcBv8nnV
LCKdQt/x47ZhT9qXrE3QQdKOmV81SRtiobgb4Snj6ghE5CusuJvd93zaG2WB403TPF6ECflK86FN
AnYrZQv4iv0NUHnAt+cW2Fq7E/AEYLWd4Ejv5+szxcrMvDBj23k7W0eN6peidurPitUx/oZUczFJ
0dRRrHRrpyU0sX4korHTzqh/gIrL/M3wef9RfR77R/40Kv4Q3tgFTD6/kns1lW+sGEKoC4wQzLzO
1zIZCFWbIApcnYDBNnZMFQ7j8kE2eiXlg/lNnKmdmUvo6tfWFE0FFcc23VlnnjQMphrNeDHz/P9g
6x2pRpWkFvlhREuKcgx9RpVxH96UOX/f5tkvEcEsTVd/KsJ8Bl/acGNFgcm/DsFTKuxftkuaa7w7
GXV1EO0dc5/kByaU4vJtsD/72hw7AdRkzACnc3LRBk9uY8Dj3UrsslykoUx5zQVGvjxCkFNGgasI
NoVQyAQh8zTLC1yKqOncvaKqmc+uGU80mm8yFpYyrPN2E/sGJX+RRZB8M2tezPgt4ZotY4jquxQ1
EvUrhfQUsT/+W+S4gqSzyivNCnjIHdOu0dN4UJgJBDolQJXz4i7jk5GQG+C1lTdw/kX9QGmqQ8n6
lzYC3ALjBvAd9TXkXSSseCPKJukK084hzgC6C/gNUEVHbsn+ZnGPUd82cs/h2dnvYcWNKrILE1Se
58dCGhMFleu3YUskDnzkSEyII1Br+QuSo1ZfkyTxlCztxHaWS+voe1K6x54EpjQ7xxfS+ovYlRLB
MXVh6sVU8qOloGRUkPZbW2+lHnwJBOsC1BtxBhUsTc6ddXEobGfAL9BVObEii+sgR4qn2h0gqkGs
7+J+CWKs5KXrWyIAwzUYZEpjiMEH4+oKNqzM83x7vuwAENC7iLkWjhDrKsDn4OTO0eETj2Aw2R8K
yWbQkPDKkOcVdPbB0JOisjYE/8+seHL8eRroQ8TCQkExoYZBySHiN0bFUQoKwxZGZlm+p2GCRzkH
Tmj5ULaBbSOp+2DmO7L0J9vSxsu3c/SrQD/o5Ms3yCuUVB0Iu2tsaGCrm2s/RS5K6U9cvzXJGda6
mYIPZy9nqc2tDBsD0RLNrzxPKLussO4YAzdCbMubJP6C2gzZmvuPSMHAHDSMA6wgEKGWMrWIGwbH
firYDG+tOEEigvWDe2Z9sPDvz2U4ZQ/gBVxM5rRcfmidTlBGeqib6zQ4ld2sIe9/Cq/XBMfD5BBB
1paoayaXUF1qSxDzmvSgIpZXVYZWYRZSEugNLGtWIy85fVVpVqIBuFIDCaukE4NsHJzJQ910eKoU
00gpDrwhUO11LuM7vakCg0XeH/A8grc7Js9rZMxf+g5HMZV/el71Fr9YOmO75jSbOKWDBYSxOxvb
b3hELfGx5prePJbfsrwh4aF27VxPcn4ocmGIdrUWo/MvGZRlSVvbvieN4kaMs1OzjB1WielzBlfE
KDSmniNRlqWOiGRQfiLvW89dMGEOnC4iqrE+Jk0EloN9RoIfTyaq04AT15ktKg8gYfLVYPWwo6gy
Vv9nwOwNcVcl22lzT/I59B1vk6r1/bggBuTbArSCC/9ZUACm9OUn0CymtY3lC5TMtO+OSYBK/MeM
KB7jFzQzjD29Fd8PL3yISfVb6+9P8I7+C+Tv1Ft0Br9sxHORsdQC1nQy5vL/zy9MJP2463OCzgWJ
o/gi5fPmshmVIY30dniRIp4ElUVbtaLHS0q3H+fyatYHb8AFexxHDGkYmPrFEyb0g7aijSnLjGYH
FwGhmfwUZ/DRlHtrdaYdxiB7Bb3HVNbWripv60o6eXr4HwDgM8ynbfCgKIiA+UrhvI7H2U4h53xN
WUBke2ESPpueiMOJcIbcLV1ABcbCJe6vHa9FCQb+E+FxzWYL3iNK65aS5FnrlZb5RzXoLM9wPxdr
UcRr/iM845Ucg4HU9MHPy4Y9pDZy/ZerHg+SgBD06urbE0B6mef61qVRS9nayLtY+ffXCnK4djva
9j2G/4Zx/47WA51da93i8OvVPBC9CMjEAO2sVXJZezq5s9iiqWDZTmEBdREI48iYo4xaEj7tCL7Z
h454en2XCaLscnsvv2aBWcatbuqdRVjhGE5TrbarX6WO8JKLfrvtm1PLcQN3cBhfr1Jokzq+HkEN
73eSSguetTcY17E8HU2UuJc+QVokytugrfZA4rsyEiIlSOFR9baNK2PNVMQEraU2Au5zZ1Zu1YHT
c6n7wVCknanrxaJgvjHpf7cX89mtU/w27YcXv5yoZeQNq3K6mp0ZzKKkHzLdqoqs6qKyCwlU4i7N
kwfKPKl6DoQGHRJFuUKmVoDUlFjBrVd96fNtvtqOx+hA6MCnroUHc2SeoShNdsYjcyMBk2rDgusE
WTbtM14GAKXHGdJx0EiotZcLzxHh+oWwhJFTvOm+XTH1YPZ+wTLA6Z2G5oQNQC/aVsXh7hFotzn1
n6XxJTdX2TY8Vhpt270nwEYTuo1IRVvBYbJ3don3wioQiAGE5PfkKHOUQLrWUFkUMeOEjm5uzey1
wQUSW6G8CvEoK06jrpae1Kn79q8CR5g00ECzPUs+bNRFptsp7kbWgAqnMZVCRUn2OT4FasVTF7Va
+9G+kmiTwhJ8pB3lFmXtOWQ5EaTM3GGQG8FSmDkm+AnYxnboiGAbB44BA+ggRKH5UU0ty0uaiN2G
O18rpttf/qSwi7gW3fYUmIhn40zKm60M5FdGz+x8R/8RVPMQbiISShPRUWU4ytO+1pxK0WTIE37u
qKx9YBfWrGYOamyRnPUFrhcT0IKaYXDYwW+yHZrkjA6JH6N1O6Thqw97+9LwL9FiLmrFt+LddW+k
L9gCLcgnmuhQ5dQDG2pZXgBXWSRfA/2OcoDl4nQc8TV37aJPHJje1MZ34NtcaBiPYkr9BZgB22wQ
CifjgitThgPwry5n/aLVxH/QBVY1VQQjOvskVbzsCSdhblHNlGmj8UEz+iBYSbScQvsCHeGYsIKF
uel9TNh27VITk6xEQzIeSOiNJzyG8TL9NTbJ1rMp2pSoRsbGQAKZ49wIGtqnB1LAYO+oxavmUzBM
5RBvTJ5INax0qER7OdXFaUXdZqShTotJXK2hs6xvVGGEx/iCsx7U5jda6cqV9i10iq2uvWXkwBUy
UReLv0jU5tHK0lrnnaIUBIKPO369XJopYgtlQ77UUpijvovfj+tZcOy4JjAAgxABaxiconjupjKS
zgOsbXbAxUDZGegGGmwB8YU+mBq4Fpjo7sI7ogBTwTgF1+ldfZtCjPbVU4UnUCxJeyLkWhPGtEsY
nT+xtxK8aMoYTJDmy4BkNpfVlLz0GOdwEsmcdeBfuUGgogsE/K+DCVpOi7UlQalXTSIuzHDMLP3k
TdilU6o1JNCIo/uNwYajRD3aAyYx/veJ+TrG/meUTGhLz7FRCN+kkl7SeFJDyFlQDhh8IdPFQVt2
Y52nC+cMWlptJfQhdP3VuPD0AgmXrHY12q8JBJpazTh1t2b4VuC1VKjXmO9fVMZBUSrYokS7zD2P
O4YV6509KGyU7cno+w4jXO337Ug6HM1YKZEZ274SlQL2BHuhFmGuVPDH5k0l4LnJfCbq6hYx2BeF
dXnGoryO01jMYz0XVi3/+0yJMEu950Z5L/mTadu2zc22uLHJ2qgGT91heaYo2cdb44y3BvmRVrcN
RagVzcxskLxaKuNKlZhRLjxRgRoMPAxAvRYey+kIX/C1N2Yd9ICOYRYqaoOTSsj+zeXB7PhQzcg7
4iJ1D0aS6gNeVYDm1LS03EVhw86+aO8tlu45Rd6EGZkCsyZvrnXrbYg8v5kz8FItQlcebJf+pQ83
Bn5JJOowb8SFcM1nDWOj+33dT9pwYMz9yllf0YvwklInMJYG6mfHEELby/mjFAgo4OLqRloV/a5s
VlH1DglOYMA7cqnA1lVvSdJq1YmILhHo9MhfMbe06/RsfWpxGrHt8+AyNtNTFMYj550NM7lOc/vc
qXbju3NcA6DKN/Qvm9GuyaFfp5QhsUdLFki64PR3CEh29/Ftqve9D5cgm2kelVTuwibqcrQ8467T
l7+gqYe7EcRUXPnk7msCJphZQEMUe0SYqRlfGcSTjNTDKkClaA02CNtoncfDxdMRxrXod+lssGMM
Ls5+HyQLUApf4zyDtZXfMhUjHaL+3x3l+TJCFvF3biIoe+W47APqlq2IlgLOp34VA2f9r1TFvnqL
SsHo6ygMwauvDSt1EBVKUkt9+4m9p07Ri+LInJAxzcVZw8H4tOkiJeQa0CshJDjJ7Ngiqv5Zi4X1
pl8kHqdaqy3tMsIsUQAVYukGipSSFBN9/faR6gw414Dg0QhrhtQjhrh5Uece+/3Bb4wPHVewKjag
+/ynLXyCC8/iA4y2mULwC2vBcJlCpyhMTSSAFJSi7pkh4K3Pq90aqZyvsQoiSL0Z34b6MmVT4fCO
rz/lcxQX7rdnPapU+oGxsXGFaroKwqchD2WCqX1ou+1hx21LyjdkJcidA5e8BYDYi42aTvzOaCND
ke+P27dviMzvWpSlOYzbHZuiLl45wS1kTsQpQDEMx3kOtg116kBsDD/W+uLENRkw0/tmcGwKB1mj
lYnxFtWfQfU4bJ22vO846FJlzOrDvZpjxKAKrA3TK/eW0gknzJXEG8M46fVpAk8SjKxSSIXfDOuv
V3wYwQlLIgazz+eWthY3bF6k3xqj7aAfobgkdSMfATrqdFRpUOLAGvHdw9oq0tsbHZsJ2kE6Tt69
YysbpSf+36+CTMF6lgUVunkqSWiEQmTPSO/ZLukH8AuDNpyA7dVm+s5EYLS5pj7T5JR56KnU9dVs
BNMsBe6u5tFCGc85xzMtDm3cWafKj/t51D5zp9rQVmfodOAxqQh/Szcc79Uh7FlrXj+AX9xuVawW
mxHxfmijmnVRCdDx3L9yhWeJ53tkNrj1aJx2vEA0AuOiEdI3THt1jSEC56V+ZMVWYKtv4j6C1LYl
mMboWS91dAEVOdn86BwGAxf7ihuHDSQsbagToTGJlfWa+bELCa3qmaXrt1NJQpuIhKBuY18knXhR
1ZT1er8r/WwPF9n1nW0b9wSU2BHC3sNwp+4zkyGVYUd1P+L0SkXaLZSnrdO0hiItn+07DlpYApjj
2kvanj/XrU5LRXUN+M27GU5RGnv+La0OhqQ+FMERIRD/UQy38Z5rAcg4M2ddXIRc/Uyps3TGH8if
sA2EtWE7kr7l0YYSJFtk5pJAJVFBk8a7AbCDz78yyMUDA9Z4i6mldi3spQcHFsO8Q/y5B4WtQuZ3
ongBcpAOkfbgGXSvCfHxWqP/vUfiXkvTuh/GmjesNEc7Ft3EuwzmwLo9Yt9bQRGRdedpHqmNN0J8
Nw4CSpyRshmrvG+aFVDAl/VuMergY6jYkFVjgbACf/50d7BQykrQoPyRvHF6hz6Wk8nKPBTdRXuI
ISt6SW0cn9ty8S6qjMz6ljBCOm97AybpTvOUI5hOlG44aYhOulYK6hD50NCrqBeF1pKIF/1BwB+g
4xayWVXRn89oyvtiNtKgYRfeeFOeIfGEbfQXA9ZYFzGcusskFubGYyrUvqfgFRtJKB/Pg69Ia5Eq
Nq2TXodtOPH9oFUpjvKCQ0yJZpjKgaBJji78HPi/J4Mf7MODDS5ATAjadrFy10JkCV8KUyksO+5C
g2obedbfLzLC/kMmo5+wr29NRZVef984Ev2vRsKE2zq+wBWR/jcS/BIaK7l4fWJbkpCfjVZmAxfc
c2gGKPsbPwa9b3UpDd3fLHB22gKXjNcrmusLqaAsTcuTuFHV+zC2/8dAbthDl1QsCKFegRUjbAjh
JO5HBoS8gg3ryCy1ioHeVX5Wvl0/7xyNTDOiEgFGc0YLlcmUzHkFE42WSflqQ0+VQkTczGRDwJM0
qf5ZGTE2mMoItjzJMIWU0sVKH6fUgJUaZ3ClrscB0/mO9cjanW6x8um5Bg9yE/9ELhIecQlkxory
DOlMcXFYRW2Voub43bLvexnbhvq8DimPjuuYGAM+lPZTc7xxctx09AYWhXKyswoB5eyRU5cit0Jl
6o8Df84ZZPJ+2hz7QDTiugiopZ2VK4Q4LhnEKHpd6/5v5r2n7ztYi8LPx8Djfos9DPRymGodyNPa
NKnda+Gpu6nUgvw4JcjeSU5a6+CZCN94umKM0JRu5lDeX+3yj2MSJppLRYIZaeN3Gv+ur9ld+Jbs
NomtEv1AfRAe/aoXKongpwwdH4TLMES/MAG+aose7NF9tNU+JsbGJZYSJL6h5rUTuyKdQNlO1JLT
pyb4CsE+BiJYRTcWWlLV9Rc4A/SKZFjeTQjxp4/s1aDhToDksy9p1jNnSw50p/8xGUrF/TLyBGrH
4cOjLTFA+xG1JhDA1Mb3u39eDJsu9hWpq5/TIA35dTOkBEB7jx2er+BVJCODBRKwrBceez8sq8TS
J4GjRYwrWZVLLKblr0MLQTX9JX305FiIS1EZ0PTcINsy98D2al2B7+fYWld6rpkdgXYZMWAuGope
o0CYhPtRu4oyH9aaL+Plp7+JuOzUFccnaveFo+xhib9Ekdrvo46lPzlheHattqvMYKGScHCrb/+2
paT0sZpuPuD/nomhLs+y/QQ+ziym1m8sEg6ayoQQ2CKsMKw3wX1JMFKB7gPTIMgJliTHifi6BTKg
uzkslIrd5Z51a5JUf3LPWuZByFmZvlQbB/NtKoOOQuT9tniBriaWP30MAuU5AJJ1uMTPEAtbe5OM
f/4mcuHYNCLdswe/GUtLR1nlVj/mcfkRHPfq1hH9II9szyK0LHQy6yXIB3qTgVNbZHLSl01O+BuZ
r/jV0NcEuQjQBXEz/ruDI8z3zyb0aJgbHF8d9LNQR1WS45VMLCyr91bVFxcuzWAQQaRAx2QfTxCo
XJhiZoo1SpHVej4nSQnQ/dSV/Rle5CnBWo/XeeSbjhPB2kzdgBDr5+hVFfsH5pV40XFXcIdNb/2w
PJF2lRb571rfjWBO5F5mvF/ohlsIfDq31LDV42gFIG2Ojhv5VakFwKzL4u7o7Xx2kP//lhCAvlv5
CvmIzHI/KySmW3+X89wgjygcWD5lcWi//Ob4y5JPwABdmsrqWNTPxpRAfHiNJvmJ6hVeqadbB9aR
PY8gC/VsxSkMR9r7aEIeacdvKL9IPhKM673DsDLONjwnlkMZBn+hgSV5biBKLNjJTKfdn9yMnXnh
M/O1nBRhpDDLjNsEn+7Hl8AyPKfC8KoH8LsmUTMt1QQJUhla8alILvUXvkskxEM3dxmID/1YTx5J
S3Gl/OpQSrvAPDI75uHl3RDU3S3Z0oeHTyfR4wMfG4CpAsfVIgJQKxdoN0DWphRfRUEYx096SUuW
9VYMIrRl90CkR7xfsqIWDhlwYeFft1Ci2ghERA/WFwQVwMZIxevdln/mXfcWnLpyL8dgpP3SosxJ
/Btowg++z33erAuqST31mNev7DPBpILk2BzXz66StkPmNSaFEnKl8LD5ZyNImqXEW6+FyT15xheC
pyi408snnYzbZUs2lw2vLU9cquCrkRGpgw7mWHrIWRdtaZXO80Dzw1FyDBHCcpq4M3V774wEcCa1
6B2UjTq0oBbmlCNbhJR4f2mDJakpUpZGWxY+u0uac55RZeDEX7s48F+EXOCSFgefU4bGIzdyTBAi
ORKxdGC7iT3o40IbQdwblYst2/kJ7fWDu5J5b4TK46X5Afj/aG4FaUoiEnI9d/6ATgTdhxjdrMtW
BlBxcwIFx3+3zVI9xgg9eqrcKm9Wa1fTTOqyNW27jMLosVk5VqrCNiUpDnMDlzKu+/QxFzeGPKZ6
pJe1yFDyYNSA2BxTwrOWhXPqd/FN86NOtMhgiMpezYjTXjfmsK9DJXGuW5ltiAfC+3GX7nnj+knv
Ys+nKeyKHh7kFsUJ8W0xyt4We5IPAyzeyrnGjWhIeOMfyYmtMrfmNKjVmbeLz8tLli5gRgvUJjbN
8ZUoaTUVuJGBafG6VRQmhFa+KVUVcMfS19WW3GJwAGqdYcOtPAlLkUa/53pHBCfYbCvfy1an7737
8zI2TyDNTVWVWFKYo2wg0uvs/X4gtuGZl5cfaJTeVbdEDkRj8Rwa9Xks7HAHBK0nSUv1G2Q2tIV3
fn0OIYpOwP3hEm1sIt82FBZ1FYu1X1Ex/gtfRELLqHe8rju54lgalFFg0V5Z9uByi2BxcdmE3gvK
1qoFUt1nrFB/J8wdr6hBBz+GfcOJgipaPPqSP5ZlFt4fD6G2Dq9tQpfenLcLbB5WeUXBs35zuy6H
UYSNEUS/eUBwOY1OKHCDtbyNKrerq18z7qmhSo2kWWwS6f1ABA8hOXT82+OwBEWnd/MTerlFrbkA
m0G+quTK4RYLvGmjZMqiXYCGYKzOl6nzdmONV6dDoqQSr4A2S37rFBvwkwmX/hZxDjp9lVejw69b
mn9aP9Csa3ZgJCJkv/aKACoH5WGzmnosHIlh7QRU18j06TNykxlTWtIEMH3rPop5dmMgtLqGiF+Y
dIqOXWzxkPoRpV+L5+0KjOJbQezdGbjiLQ9qB6Tq8VMRUtHCFhR8R3Dbc27dfrfA34e9RyTvpmWH
QbxUspYMtlVAebRFIWTL4xu4p20eVHzw8o5o6Sa/jEODXleBrQGYPTNgwyPULq700/W4GazKbVvR
NUG8IMLNRmoePODEvNRjJi4Wm0SIW8lVPb0vBajLx1ghCuCjehiCvkwLdlWcDNedK8Bnxj0OF4Nm
heo5mc/wQDO8pg8nOm2EVO5t0E2c8oVw5La3WLthoa+Qkxg87FUQDXkTETVFhyrOnsJL68EYcKfR
88u5N6apIv5LDWlWGSwh8Br+5bN4LjV2bRnvne9KLw8tjZgWsMQTPWtijwxUvtdpaLSXAidb/7ns
GH7privGueWz7URMYbSUepo3fniY1O44ewAk7upizdJaCBsyuaXH+So6ztSwzJv9f82DX5+7pMa3
EPQYShbXQlQdUtTtxM3eeDgE8c6XYYe2ejnNtWtJPdWgUKoQSZQ7ubRMcXVQDVPIN8/0DGdUWJbc
JN2oWhNPguMirkITI68KF4LokIlxtS7rGMr7gy9PLt/p8PZVuMYMp1R1wV5ngDL1K1qx26+ZMYi5
9lPIRYZPtw2OriMLHJqszfBqLXrsxz4g5coLo1/b16O77LiBz9mOQo4j8zjem9FSSDHu9Sb5E4UT
ALpkuiZdStS50S2UvJKcJ9M+YSljVkJtHYVYlBWceCilQCXrXB4yrYhAt/q73FpugxVcPXKU6ctJ
eCTTxALUfJcMwGVzuyCAJFVocQFml09Iao2cfgpwjO3mOQOGVdbRrKRyGPfYfxy54zb59dK80GOh
xBG4G6dRT2awsgmebA7RUjEtBsEUojyDw7l+8IO1rkPJLgAEKsLfzBZNnam+mc80xB7NkL5f/Ec+
EMsgrRXf4Uwmg0KyLSIOcWpY5QQuwD9shyuveZZOgbpe34eRoNjN/gIoeFW0nClbpHXsKhXCfEG6
IiwMDdtV9DkjMV7FaZw9WkAIxeLHFrKxVL3MbIYmT/8a1fj+fLyKejxjR+IaFOtxwYBUrCFpU/zI
R7qRFZVbjlMWSZilg2LkGrLCHL5ae2YK3239dwkpgma2V+tmKbkm5QCg3koTUpMao5iAqdVPfYGX
KXeDu/2ZAzvVmiGCUfcooxxTxZAQWJhxc8P7yGCY8g+XU8bCFRC4FzbjjBC6M7QN2OZQyOlSrxsI
8b811MqLztHV/FHRRoVKukDOc7dgyYBEzstEojn7qBOJyfNBlt86YpYrayddGSWXi4ogkubBVbK4
NSJi9HMw2aiUnbyeYwhXS5oTzggr44fTGfv/6NsjCXIc22Nd7775XQ3hKdf7NfCH5dCmb7J+wc5D
j2VpKE+RJibWu84cVTKz6JfPxldxfm+DHr7AMsD6nrTXYEEbYThlDBdWtXIIrOlzU46LP5z62hIv
HjaMCcJEyroCbltUaw88aeiLx/gsODoVai9m6/JTO9lacZkBQ/VL0j4Rj8jkLqh4/nFEE51fgaap
LjDkvQYZmCuCogDjqBVPli1lqCJjKl/k83PAiEDIycd+TgJ89e607OihJIJoN3zWCFGcUdaHEpiK
bqkOsEvucDOdQuUcxDQdu7t1a/3Gm9iNdHx28djB2XInLcm4QeqMSwTGbYDRGjSWVz0CbvGGM0Mk
gJGZSqQWQnu2fQKlZ7sBM6Tkan4rBl+dxU01l6O4IrZvd5ZLo/avuazTs6ezXPwmDE9Z7Q0bZSUw
M62IKg9FsL6xD6yQLIya+ANoRCm9yyrshBSixu/VLWzygIIRtChzrUDtALc1BfLtnPzjw/z7BmKQ
/0dEIzxfsTfpWznwt/jaQlAL6b2Ehs163GOcJrFY6kiDYIV5PrmITDtzjqXbr7NWQJ9gerrFTA1N
B5r37kXU+yZSc56FQhMgFrOc3ah8ynAqTFTPODJ6YqGPjqhx8y1CDbxpEx4wWGpuPnrDltahEj89
gGAwQ4DadbrKKBR2A5MoXpO+vnrVN6LlglbdyEtch0E1AKdTd9N1tjpU28jozWpOR603I1PLw9CB
Vp2cw+mgeT/5qvFxos5gQJvXjNsUwsxAZmR6OM6os1nUztn9uPt8yWyhchDFIajgbzb8kC7eE51n
JoYdDG9/nwCKishjy3ke331g6l1DpluC7LCEmKp3SMNcEKs8haj6QQuAnPoIhLAczeCb9xCEMBuA
vBMWtQ04paca3Nho5psRf3QKDaT78C+FKbgdsXp6r1I0rPIZju51ZHmz+70W7a+mekkHJTYBvZN4
5a456oTm18Z7gm/bs9udCMa85QMbi82p2PXXSx048WDsjssJyf5CrjD8bGX8FcqcA49B8gdtICBF
A6tOPVz/Uy3sHBEoxtWT2VaUrgC3cpEL3xoLEbybnBSOBRF5PKT2Agc5f5kgiGDQJWk8jGo2shwn
Z+PREgtC1pBaED2lvqj+VwF+fKY59QDZZ5usIQytBETGReAdevxQivv+n8lysp/9c2cFO1VUeNIF
rsRCFhhFN+KdYq/S49sKsmJyWjv7HsFxdf9p9/uB2kKRa6Zzh4EEaDPEXuFD5rrcFmhZYixEBDjE
aa5pfkDFy+AEFmgLsC0o4M69bFeqpaHRv0gZ8uB0/gTZBdqCOabViXQj57NGNJhLA3bkP2v4eux/
q0lHo6OKcXlN+8pecz7X5feGC+3AWVpzFuvpqKk5x31/9JPhPqOuOSDR75gewmNQjAIgj/ukgNx6
R3BdS9iN8jiC6UZpM9h5DCARyzXKlgeXVTvlTp79UxttCygYDVYuBeKq7aWIkKYy23MBNTz7AvPR
K1yZ6VYg/W7aO37kmk76kDI0kjew40L1UFzLNGyzkWmNzd1INde2zX5gBUVeR6AK/BfDgC0TnTLO
Dv17PEJHJ0hCfhh8GRyhnmymCmHg+FA9AZHxexNN210TBf91WQS54BV4F8Di9gFXoJ7thNwKgNDr
RmcbLadUPyprczGslSsNigzySeSqDHCzdR1fhYsJVIUl0mFfWD3uKej0nUpEtxsvJH7lzUVvmfnQ
G9vBUuSsue6ZT3PuDdQVCzqwhzRSdVcd3/SXMw5xjL7XwUwVQdRl3rBowkS2sQH0mc6EbI8f9kUl
t0qKSDT7Fx/j89DBqqz1yMyvF/dX+q9qXKb8DSF+X1yMQgdSGogwb5/IEZhDPJGMlATrB898f6bA
P8MQibUqQrHQJvVYQJUdTbmYc2t4qeYuOae59fq/nD/EgbK/uxbKbMo3IdJGwQ38fzX6bdrRjx9T
sLZriAr2rEphcpZpvrli8LpJlIoU2CMkxLwRr/a3IhbcDwtv1JptqgPLkopAGb8J7i+yGdXB/kbk
uHNN8wg0yDm0NtUV6Y6EDj0YvGe2xboXg+Nza8PlpidKChd1glnn4Oc7wpb5G5VNbO+HATrwpxph
GGP1Iy/4DniwJNrSfQcQY0SpPTa9KBgFQSNrCb2eRACXPYyY3K68RkHTwuk4mggQdJoKb3YNk7kh
C4+Cia5HH3V3m2PdU6IWAOjsnWz4PF91FOAoAx6Ng/66lU2cbCUUYN9Xh3pyvfTwXuklqVSz9RfM
qcqeIDxQhQjJy6i8U5VRIMwKJHq4IF0ktfZvjSjdbHV9/MSQjThRmzrrafI016kdmdAmmk1ILiTI
02IQeHoRBrS5hQjo75tJyFae1tmffAJTdWngXHs6qZA7z8duRMRNW322p6jOkCJZgO4sh2JB69sU
t/guwOzKIR6NVHPmwVzIHAOgMP/8i3ts/Jmy05aMaUbodelZKhgPCXZ1xLANcfIoWhePfsb6tGWF
do06xqeRBi3J4ieb5Fw+2fNmvAAL5z9rahJS6YzencHzk9gacF3ZOzlWiIp7b9LI6DEjdv/SfEn2
EsHA14FXo9S4KG7sz085ZpYiASVGRJcN5OfKsvjYRg/czpX05qpPRXA/EoQ/dAsqTmoDaPV/G24m
ueAfivcZXzR906h/2Q/gBgjZnEQcmfDtncoFdvsRZfNRP+p0uXNWbbz1oPFKVavU8TbKioQDGX2e
BImHxFNlfrcqMdBCB5AqGMhfJ1PA+esNNbYHzKxSpxgWHje/PvolJbez1ytvORaVFx4a0Z9Btmrh
AEBXa/nwliz8oQ+BwTIpDSoJtblaRnXQjf3inBu5cZi7Ec1SFgc8f64VdG52sdIANc7rQJeTOQqF
/uR3N1/L+2/vkR2dB6ohf7gchBSN7GVCvAl4Qmu0LrmUWqMRlq8hWZS+upr+UFC5OD40AfQ+tePs
YOs8SA+8Kf2xOaZdU5t8cripSqfXl6qiBFl6+7Qz9oDjfSIG6VUrlHiIzZfCJTKmq/KfhM+4A8Vr
gNuEXKi/cMbOr/BgmRpgOMEpn7NW2MKpQcQt4bnFIrDRkF1/4AOJwHmIax/QIHqmiJAjnGgZaqwD
sbYMZFnkRt3Kued4bEHN0zPgdYOTKRte+3vXQcQKBLpnslW+fV052l8sn8EqsFAegkfVJ9VgAUo3
XrNqBP7BnvMxYGGlMvxG5dVM2ozX/4X4eJcoCsP3gCtnBmrF1tK4nOdw+q3WNG6ICXCkH8CoEwRr
U5k912lCa85fDF4VMSrcT+YqA6A8L2T+hRVe+89KyVWL5i1NE9yxRitywvUOB9+kBeIeZLFBidha
cOssMk6lI1Z03srpWEdd6jwcxPp1mrNBREwZ1ze9dX6nLSgVjBNyhEF4OLetu5SMu4vT1fvtGqwd
9UrKnzxFeUD4Wc1eQ0+2TxIlk1Stu2k++9E7WsWEQmhfBqpbalUbwepFWMFtyegsMhxvT8LjVVJg
EWf4JC0M7ShDnYHwm+2QAwYYvLQeJ9mHLdzrGmPfpbYgk+LThdmKZEMsX0TtQASCZwweFMWN9PoR
c3SERAjXbBGrwMpyc1zSfxI8vxhItdXWsMU8NXLGkqKXOK8miauIz24NJY/oEokOEKIP2WzKAMSY
gqThzViiDDfAgam1Su2iemQwBZjgNV5McGA6vBNyXy+3JKfU2Mz8o7gM7twI8sdtZ68EiKMYgmnY
cYut4vZU2WR5epvAfC3M/pw7kR1gqSancJSNP35eSmzZ7B6cefhEL0Y9ZZAJlnh9+FPBrbd+fjkG
/eW28D7MBbKnfSNrUvTAxXuH/8SYvXF2GaazeVloqat+RgKVMMqEEJDKGF7jDrVbBC1jAitpInf/
bhROzObS+V+6YAJgqZ2+ArtiVHeQoYZqEwUU5nQ5IYoit7zRO0E8fclw/W8loG4A72t532GdjYa9
LGgVogwl6hBQ4SRWC6V0LL62WGk/8FzNE4H//OOrjgS1paRzOdeqcux6eEFsOjGyuyQnIHKIhn8H
u6SIw9z4L5sV5H1FfMdKLbOgEuGqhCYJoJ29BISxVfGQzKVv7QIcJEau6td1VrrpxSRWthcu6K2H
X34vMQcRm+znoVC2GIqN2TzlV/iWxNhIM6uQT0sfNL8Ftuo1L9LkSiWYwktEs5cXAlGnDCbUF+fg
T62WIIS3CXCgbpAyoLR7Do4VsTOdMLvfZz6zfnNy0XO/KJyk/pyk5V/ADryENQ3Z/NB74As8w/2k
TfGxUNV0N92LFX3b1Hs6N4BAHsYaKuiDslX4D8ikD66alkX1YK3GN8gbEmzsBlQ3KgewDvKw4IEO
PLsFKNvgFxcquBh65XWmN/6qqQgHmb+PqcmtmGbBie13Oidsr8tHjmQTaBNNSJ2UI4m/KemQL5TR
/BF35R/MNLwh9G2Z+593v/arE+ZXZEeU4lXET6Ai/IRoIB8fMEACJ3Og7UJSng055k/zQzCw3G8D
icuAtwbZPidRTzcDlLZd0Qv+3MbKgIEOG7U7k6hYbLlqGcjVhlwVNCc26dA6CqeMrNcpV76blL4D
Qmiec8Qz/dxVl5rN4R3nglk3gtbv8N0TaG6BCVZL3H9LIxA3Q1wCnRG5MKZn2RFC2jHMKuJOCzkA
IQiPeDJZQ+a1U9GvjWW8OM5bmzIsPclVjCfi1060Tkh+GsOEpXeUGre8O+3s38ZCORkzTT6wbwP/
qtK9+nRzrBTRsCgJhBX05BavU63jLcL67FND1DaIvHU0GxP5Bk6g7QSkAp7xwlep65ihkhUQHRoO
x5fV/nm3PetPilnGydgLZFvaTYg6T3H/ciwN1SZKSpg/MUo9v0slX64yyOlfZ2t1+oMRYshUmQfn
s/nZMbGQOQoKx0/0Oshov2bnUZZT60LCt6DFmCRl7GAyQIOCZkCwpn1UqIi87ilZFl3anEuVYMZO
VMTuGQoOdZKjYb0kuOtuYxbO03yo9RaVgCqW9OONe6a2qMROjHOONgmU2wVi/pHuKpoayZBf1CWh
2T8pmdmfp/m8tj8xSyuVqKnFJxlWWDbhmbfjvbunRU6wJKFfM2D3UNCiTs6xUBai998ajXY/HHnx
1yWMPkztGxTTJCySCxdhqiB8SgFptRWwhot0/pbuogXrxVKPViRA1w0LBilpJ+s4PU/bJ7+cLpjU
yQXnhgvzjouL/UD1DP/DYzNhrBZQb6XUMcz+WP6i8GzOsNCF/TKdWa3P9OuNmJm/YJyEQPzbYsw9
LW7vXC4B54nT1ow38uhKW9lLbnbMi4lKGl8eY02rvMeULB6QxoJKruBioEJjC4rlQK8mRSHvRyQi
iPVf8WR8ChksD7WdW9HthymaUXHqIz30PUZGfLGSjvtWyXdZyj4YQEiemJWbf9BJiyjVGtDqAzOn
KSP4MLZmUvl+Dkr+7to+mkmBiKG0Un7187CpkBRC+RMuI/sTzYcj9zbrZIIHsXQh+7YEH2W3w7N9
UJS1o+EOZ/9fRL2G7Wsuc64Ly8W54wITphO+gnaPvphFIerBFezqy38sKq/oZh17M0fFaqHZOuVl
9116tcEMaCsU68KNhp8irkZvXpZNmIi2m0A8djMEdKd2Qj/E5DSXxJetUAXaS+u7Oq5hd8MvtG6h
rD2aPjan5QvdceWAqf6RyyRPoY2JK4FsYYQ+Mh6v6DijaiiNEgPrmTSnC3XcDzFUFa6UAdX+TPGC
eYpaPHKDlnWIL1uMDYnXFA8MwUIT1CbJ+bDEY9XLn4aQIJ2aaFbjDQ1c4q3AAWHUnIXmdmtvSY1J
zCOY1Y53f7eTnThim4EG+cKC6nH/16x5/iVLkRrAsWBSm5OhxuRO4l0MrqEeGgM3UoeavCLf7F/o
yqMxTK8eLIRL32W2yEOrk8LTlwdqs1b+jUCyqQawGJ5DzN6zKhJNl7zk6sz6e1+VUDRERBYN3gW8
f8jz+VNxVy7tXXwjGA+wmUma91yfKA21jEQY/Zr1OJVNZhI60RzfoaApYemzsiaHadX+Su6XjAWF
AawM4WvXgaenCj6xDVUMLHOoj9rwmePjHWn1PmJazg5i9PhRG1f2SlzmiwQmLVcSf7dPoeUssXc1
VosfDD0eaqhnO5GMf5XldTtwKlv1APvQCB5xySJe4ho2LFQm7CHoqScUeRW8sJ1321q08rDICAPr
GE5IYWqiUOUQ1xCiYviR9Ox50X3j88Ahm/YoHg76ADWmbeJuYW91yLsJh/bRMQOU/uY8q6hsZFD9
G/g++H6R0dmWKdCXaN8XPET1nNZ+dOpKDN+d3OnBqJqWpx1uptIqZMf2ObGUM0+GBiYlUa+5CLIo
+YrrM+K7l9K/NtCH/kygFnD43t6Sd09vtE8SVxZHoZSDRc5t7uGgcpKU1ze7jL+0NhRT0hweF68c
gZ5ga6yjdRdt5Dpc+1l9NTSwBm+8rTm/nK6xNSaBiDaHNCHZEFktNauB2jCBQ63r7R4q15wA6qtu
OPrHMWkVVOeuv6M6XisKFuaTR6fUVOx5f6sWFQXtMg6tIBS5Bqd5g8zcqFAhXWNE38J8Kgh+eU0j
r1e93EaE0zX4/rJ7otbNxg+s+uPO337hF3yDJiEMEwqQT8JI1BjDuSVD7fUrvnRPng2GqmMmmWcu
nADZ3fIZAGR33pqj4EOELn/+Hkcp+3cqGXzz6imkedBAZJtrNM2vujk8J7OMDjOPMlebWpnYcmTW
8RaTtRidHBoXQof3huzV96zkeO+2t7eO//uMhqwTar+VKpfzp9of8xcJaPURQ8/fpcMM1l45dVuK
uL4oLokGfj+f1v0Kqi9NoBgABqvpyzkCSZkBtIv+9FI+PCA2JIdk+rQMN75dGAnTxZuq4e00ESXA
XY9l5uoAv/rkpTTBUXU7YJXQNA47gf+vSDkKlKbsX81JJvyThx86Jj1JJ7NGV38YU5dZMMFbm4jE
tA+Z7PT7TctRaKOeN2kOUSgqYG0mR380d4AxWt4ksM9ruujhYNlpdPwjGpIXjSUuhdyk7dFnF0Es
KkJjGRDNPo4qlHp+7ILy0c3GcF85a2/7GL9JPHsokubS6CxxBMcB6UcXVgF2YRf3Z4sMl1PhauNa
HFtjPYOj+NViwuqK4y3tpTUM7a/cc4zxWazImYJktjL24TT7Wg7Hhrzmq5fbtroSCSBF43BJ5fJU
x9ziOUgeCiFzSju3MQ+crhGflAu6aP25EHwjnGLeMyTq5Hf6E/reyuAlDy34mRv1quGMmzefC+9W
9HLq7cuKbrKGqD/pTwik9Z2G/csn+Gv/nBI4SM/TRe6ssXGYRRJa+6U2w1WXIRqNpeoSuKZ4EErv
x9hTtVJnDCs8nrEzOZ6qiqg6YomGFIDZzH+fIz9NZiBNgPbe8yb61Ex4RDfxw+vmR2e9qT8Are1s
owCJ3rLPfKkqzTCerlSDkOW6d9nBpwCoQSTYJjnkLMD6UlBa7eMzwKuOdbJVqOTfwzxMzP2ID7Kw
Na+VvJz615iVbGHM3WEtFiwS4ClIhU8Rv22RvjsGAEbeFCCfaVRKbcGMMXhp6b8neXiWhzkMvvGW
N7ytX3wUVLaamKjY0K16RYLtB31sRAgrQaaIFarkf87cr/NI4ZIadKBCDLSG649rCbLQpXeyeODU
5YCK1+zz1dKc796UK8cl3k2vvu4+/XwqiFiBjhmBP3t4sX8uXeOzSySbW+KvXKLAMunqE9RuNi2e
7XplPXxp61XGvgtq/SVXu/YpfH7PYbjORrW7YCIqwCz4+WGEkCnl7ICsS6jPIbENcvhRztTjyPX2
vbmLwfDUIJJ3cuEQ7HohLJQkGGsAxp4hBS1aZ8DAWWBF0rwYyLWLsJWWE6pccOmS7F7Cquy6eOkN
PQiqzZj4DqRgvWCcgBpXuIR9D4utyaZndpoBDfRPdlt/MNE3CjsqyS6MSfdfd9rBnEH8jgeIPl7R
pc5YSLts9BzctHQDjqxJvfxE50nwaX6jaDpcQpTESIfWLMWP/avivReobtWO0bO5dApdJ4pHsFvj
WwTMV7nkSYM55yjxPINrM0EghJ25o66iyHvxOfzZutBKq+KXQ6TKjEUhwpOdeo26QY9EVhIEt0p7
R8MkH0/GjX/v/jF1XRvU9dIzvEjZXb/TkKS4LsPL9lJcl1BXXjXjU75Fs2L14u2BtxGzTyRdduIs
L9RB+5dm63lJDohdt/s1t8RsInzb6ugIPfnuqwiFx6E3J/4hYJDB6XZP4zJD/ltI/y9+xR8GZML7
tUtf+eEWyWeRCfmOTJzUXCNn97OfkJC8faVyyCgmPNwyRecmjnT01WS5scougwlpuQPAiJrieEAz
edjc7LRiGDdbqN1dF9AQr7+DuC9pNZR0uMYZEc5xZAVrRcXFftbw9Igp7kWK16BJxaGRRHF7QDue
CZJrIHAMPEqOU+Cf+mYik/sUkfOvX2jWOQxwj96JkIpfqx6sDDZZbYE3xv95B5sNQLjfId+uye2W
K3LZ1OlMLgOAJeC+mGm0rOnJFdpIQ4f+xfNcW5vx1YSjL4gKXEVqD3eXPGiW5FbIEGEWwwfs0t6X
fmPxz83yU3ysvgMjSgNsTBKkItq3uVDCzaI73pSmyf2d1P/3TUXJFojIcY6vy+DB86F7WpHNIENA
iqBZxVMv+n6BmhgNQXaNJnx6kH8+B1+Nqqg6nhLIWn/Ewq32clZwUFd8gEaPUvO7qKHo3jCsOebT
D7yafG4FBy2KFHNvpway+sDnDAt1DoL0PP1QKH4CGqGJag9sLHxzux2d5H5ez8ctEIQ7ojd/Juyb
z7apvpPG5cAubAEz2GRc3dcHhvgQPs2/LtAH4EDPYkkh8J73gzfX7VtXQPCNo8PROa6ft66Gt5sr
JQaHClmCmRYS87ktFqp8QDyfYLmjGOo1YjW19dgDRqmBaBqf2Sy4Z8WaAQxwylID12slska9DPmd
HY3u4B/xrIAUkYeayX3vhQ2n6LMr2RRDxNAmZBJ6EdeyPomUp+EqZqlxH9g53KiCLn3L44Nv6Ras
AtRVJp0/SwMQobQKbbb7+T2hHb3G49H8CkAPLTqMODStmuBXVObJsXISr29EhI3Qk1UnB2LZFGoQ
ZslNfbO+oQsdLoJ3h+00uAEIpcokPkxCJEioxYJEECwAsj9al58Ki8VJfK48jAcXGRQwHywBHDbb
v8kcwVDxMx89vftILcQFDKdPq7ygb4sChiRki7lw9P97z88TOkCZPT9PgjtFt0D5Qvo7udmnK1oW
S5PAKu1kJH8ia7Oiw8whCaUdPo71teg2+S0rif9LK8/8Y15qac9v8Tqa/3WoBdksltKd6Hl0rSxb
LrKm+6HcxvSLm/WNOBf/I6qDC3XuZvwGWChKbpFsK+cGu2/0YZ51kWWqFmEGBwvk717pKaWuLGQa
eNiGBQ3Z+02W1JYtlIDQB4svWJuItwdhxmDrviuLWwzhRxi/u3NJsusHh45bUiy3LQffl3iCFsme
rrVCsG87IKlZb6jEWkLFXPFOwnd14hPZyH4DoTtrEUWlOcCskRMJfjX4lmLLndP+UAKiHQK7nASU
/X5vhtWj8j2pd7HkqFSpt8LG/ItO0zg5aBlAROpfamR88nXaQ3VOjmvlMJRkIbDGf9P9po6haAG1
nvPEHa+tEhWRoz1l6NjPGtEY+SWMOvqAbf4tYynSEDRxUR/e6AKpfBqQxLrqLFERCdyesgaKB9DK
O//5s3lONfACHeyhLsKW7uYYoc5W/Zxvrdms1zbg5YNgpBHULrHR3ikZ/AFoSSCR00ky8Dnxn/Lo
v+OU+aB7Sy4iX2KsVJhwK0HpyXSHBUd+a+19Bf+I1A1sGKfVlg84x0ElSnmqhqsfiSSw6KEGBeA+
wwhOkZo5A88qPVMqnwjhCcX40eBoVprJZ7Eo+eAlmr79R51+wF5zDIkDj3+8pLUSbhzIZ+hepiwJ
HWd983MPM/8WHiYkiUbiF4FHQWd7Jk0G2nFpWT4ZGmX3Q4n+h20qKemqAzvOtlV0mjNrBPYQywf1
xKz8OMuMyoUbIX3jydjidHcfcdRQz5hiAciSFaI138y2hwBVuEkFV9USszvUgsKYm8El9Rgl0VqX
p/Gv2esaOr8uofTUDG6QKj2AULthUWIt3l8nKosGmDqkv5QH2GkHDqSL29PjRbt+VPlQOEOK6GxB
QHdwYILSLLnytF7ZgKLt8UYARuk1HaBjxm8NZblcKzhEdzj37modZn27BCyDhBMtCiwQJA3Tvps3
mEVmvsQmKHBASa9+8yBb9FlkS+vNV69V1seE11rKIiZguaXjsQ6lg3s/Dg9MtLrX0l7VYgLjehw0
Brnrk/2JrHYo8y59/Aa2HgBR5qVew6C2tw51EwaWG0l+/TGrnaNoBTNo14NyqGCZhclpEbsNgIVj
4/x8zX7sfw5FupLzUWH0E1Hdu8JNPrLZeumBe7I+2JbQPDiJ2CBeBdiz71sWT/FY13DDWreZJrIk
tvYP+4AfY9pW3fbd57jO4iTjp5festeyL2Fc2xOygiCD1WmZA0BK6oWs8eNe40DOz68/RSag3BoD
9FU4mtt5nqr7j69fcJb2Cen9MrTUGJlqiDNIQsNqISLaRYQcISGWSSrORGXXkaEAHQ7thaVqGBqm
NkK7grfK2dgK2dXaomFVIssBkfmmwgQ194KSajAKS+2pCtjHT3A2LS3ISoDHb3UsdtJEEIkxYCSf
bzDAqm6ywXfJQzPXAp8OSwf9PsXqvg1BmT+83fMqM31X5OWEM4xIA3+aAVSmAAS/WHKqTZINxUdM
wIryCP8a1lusw5AIuL2LLfGNZqE04cQoQKIFr2wcRtNzk0XRr02VGCnCLRX9dOypRZQuXU0qe2r4
93Zm32EKK+7E/ZF/wejaIpQf/Rb8aMTKWPgzWZ7KcxHPzVLHzuXKwGMmLUAPhTWXcJflt2Fe3A0e
klaW1T35ijn6mehPl3fMiPmWU7/WonNiYb1DXuTEQxgZskujhdyP0m0ENqq10gYfoco8cEHg18vB
HiXyr38MEgKRHLPo7SaSXFcQUwMWi1QBJw/bugmJqSUbMrLIowZ48pgaiMk8/JGABEbK+tv15RNB
WimM1b4Xxd7Q9s8deQDfHc9c3DQ0tJkES0lkwQ2EAJ2NpCskhLuxZtJXzQ+JGuVPz0HBjA9kEdmd
EOnmgzevfU5JBkEhWBeZyOzDLATMyW/sixBtey5mtch1tTIJcp4TVCWaQkBpZOUkQudpoQD/COwX
NCRgKkkpFcduc64NDSho7SdS4iXX74uPo5mjU5sN2VSSMPVcf2F96kFwS8ja+2XkRvHzuOrAQaR1
GV9dRjlxhtfmTzkGV4Nd0YxwwQTWyAWSUvLE7l6RwLaboEKRgcyuJYZe4svooCS0ZvDNPJgFa26r
bHDDCMgFpSdfgtbimPWbT0+cQkS5YEH83QFOR86uGJyp0TJG6RW02zSM6njoG5G4XLVo00dlauMF
Q/aZBb+JvCE0JAL2Bxz8IWEk+GvJ2tIpzQVkYo1hBN2M50pd4HnnAwXD7tYYtO+DDPpXmF7qPYh0
FP8ffT9qSp937//HxSMyOZtT+QuZCxIHLP/QxRCObVjXtF8BcIoqf5TXdhz4ivrTldWkVXnJJqSA
KxZOl0SY1X2WrYwsqV0cXAAacUB8al1PLbTRxge67cHaIhHAHd3JsdpdX9oGJma+zPBStykB3O5N
r1t50E85/goSU6HIaSLxb7V3H39HJNhngGrQirHSMpBcpAZJbWU5N5Uc1as9Rg5c/yHmxdLVvH8L
avyanbuhtg+l5ZAYkEF9ph5dQYYY6OgSWf8LcpUFcKH+qhqitL9TIwCJ/8hBKDPrXputngm7xqbm
tySAZQ6G14OE1/BtdNK7qmkbzqVjIYMQF6I5Mfe0YWYsh2LfsSd58Ikll/HUSixCU9HUbUz40Jj3
B3wvwLOefnCCD6lHM/CT6UH9bhlwFEP/IsRUlDaEzzeuC15m2QfT9F9rs+vAxNCxkczarInBv0M3
CcxJp15LwxER2b9og1xYRSC4TWgNoZON933Q7u1vV9/xw+rvHyZnmSHhumwZBgff2VZSpcOzHj1z
v/o/KXWEY30qHY0UydB24cP62M1j55WcF0nSN/zIasIafwGYRKnd9CJiJ7hXnBuMDXjQAC5Qa/Vn
PwlLtXBNuYwklQCbfVBsslr2YlooDL3u7rg3jBzFZDkVoyQiRg0CWwsv74nwBRfZgwwgizOIsBy8
EBJmW3YULnR569aVV4YkoGuz9JGny9Hsb0nKin6NrovbXj8Nb5rb4q1XA/riact3i/DO4lKbHyzF
pM3soy4x+XvWDfHxKAy1sM4V6yLb7dduW2t1Rb4yxpo/BpOJharW3m4AblgoYJCoGS/HYvgsuVYt
Cx39iOx72f7EXfL19+lHLNWlR6Ou+DbnuEv2wWt6RVGju0eszIYPnszujsCP4R5ooQQlyFLZ5Cm8
1ebeVtXGSm/Duc5EscrSJTRfcnjGwV6mT95EnldlYqm1S2Sr5pnFlhQNFGSXf7ZtdxBIuQS1ayyE
iEcR7ClMwh/fCtmRz7B2jZvpCx+nJ3Ta6AYW4OgA16efoivDmJhY2Vyaj3n+VWPDgZKr+/KA2ice
3J2Ekwm3CJiv/SoXhr2EtM5PB2jPWoXN9s/3mp60ANeQEIsLRX7qsUcSlpoIydbnIZANKUxELCjL
FeQB5HiljRuLBizHRIA7Z5B5f5lBNkZhuiM/5rQ6uW5VgJgLwfuzN29Hye3mB56JXUP9cfq5tMb5
z7SFCMWqFehFZl3sPXGxdXr4y99UICnVHykXlfgT/2U/OaGpbiBYtbSxaJ0uguMxVUAdwZIKjsqX
jHGkZdA1+lWhz+QLO3yEluBAyFn0nb19RPwFKj0HqgABxEbPOCqDBagfLQocomsIIwyxXwST8cQe
D7xrEMtyDinfZ3w9M4JV61+2Ogq5mWkSlPDVD68vzjycBPmFHSXe9KgdJEFXYACJFUQTGJNqiGNJ
nu/dnSEQTscwK//HjhNxPmVlS/hGa40uYYX1DGYRnxK7orDoITmYeX1UEwyXrrqE3KSMvpH2y0vI
GqVaJbf0is30JMNWUaIGDRQnOzqqI5FKa8PvTt8OhRMvoo4/dbLvBNHTQe7YLBzmbTJDr4hRNr2D
C3si8fiJWcBXOtulRI7ydnxdDDfDmyzfIJROoSsDrMWHIsCjnXqr6PLk+eN19AmrnLJkzFGfYnN0
1k5hS6fSzFV3Usj7je1eFklYrLSJwLIoR7fxaFtbiqMa1OMTXySzXZuCsnb3eDyO7SvbK5clWsal
iaPRsmBhssk/xqtTTCYEiRpUASmPNgw30raKmJvW87VEy9hcYipLo1mwfMRZPNMpdsVLGy/+vcjS
DAJ5pA00tLyX7eTYaTnagwE4PgDerUYvxOPm3d0djCwqjnONJIMLxe6xZvcbCHrSLff6Ze/+51AL
gb5gRfQmYwiLIysY5oO+SnwQ/DYMKuxCVVHfWvFtd7flNLfoxgz5XVbUS//nsVhz/o2UpdZAkQu/
Tj5ifS0MspeJ/roKSkMCVpX8gsyJpBEsBU+n6leS1eMFbzrmgEyVNp1AQb6WlQiWIQvP82InHodr
AfUF7ydfgf9871gw+MlnzViCLqD+9vOpAnyjPGu3Sd3yL5Hrq2tKjexf53bGnHFGv0GPNB4kOSRJ
iZSn8Mk3Abgs0bYQdWR+EkNYJJkmvD+gbcJCxPshsU6jg9ZxL52+MxyiOemUwP5m2iHSOOtOSoj7
46k/k1kRiV6pA4pxWYDS348aYE1S9On3iXCprRl+OGhDd9bYZbXXOQj0vNuc5VdZHoLuUxhvj+sD
/gL4B5bAhJ+VlI6cFf8NHkcQqW322Mu8LB5UCRya0y1IdxK5VfE9CfAT89lX+2igB6pvpc57e2kW
1Li93XMJ+aw7LBpkJr5DCY0BKsmTufhXwq0zKH5ar1n26hL7BOVBjUBzo7pEFsUW0XdU4iuvX1nj
UHtXcZtJchoFLoAMNCkFtAlcldYy8D+txYvN+uAjvCQgy2UTCL12j+JiHZ2t8JXduXoeJcGVr6CG
H/RvmxvKJSnBn8WbYWDkSNNclp2IwSm8ige0jX3hCEDsSHvHLGZSFGN5bG6/bJyJSe1caXvki4Ss
yleJT5E5705w1bRtnSo02glToFEK2oGCyOq7JoZ8hRpCvZefOUD/zMFROs+IZDH9ObrYbSRwnchO
NgPl+85VEto9BHSt4UC1vPSSSV46KJnMkRy77h7DSYO7C/8Dtae4SZ5IYGa2pY/h4/pHYyY7LmhB
QA1E6q8Mn5y3J0Yc0qcHPU3xnUz5wlNlm85Oc6+6LoK15PHbTXWvzOTOYOjjIPyCSv2K0El8ppev
VylkMTZC+Y4ORrm9fJD5u+KHkXYwz55xIkfflRpbUfAf0iSznHIjbrJIVxmps7dmdLZyOjQMZ7k3
3RzDy+Xn6r5klwVLVQNV85znfX+LjrfqmU+qbjH2D8ySFwMWw6tr1Htrwm6gOgVczPYPbEuUK7E/
KxuLpzf42lLinh+YA2daJDPaqPrJExPxEMNQvq9QpanLg8mWU+lCMDtojzg9WWnAp6Hz/nfpkANm
4DYq/Qjy7MuZUQxfWPBeHLrZBdkn8b4UEBzG6aAQuvdSRpsveiSvKSD5SGkhxU6Jpz9EpJPLzKS3
lzBp7nzYHmwWmmog1ELjxyY/eV6a3BvZYOXFaQ9d+EiFymfVeU1It+iWu9UT1Pd3FFYbwM6oIwpe
l65g1U82RPsLuphyfxulJHIjhPg6xHvlBq6TonF6L7QBTmTOvP7ciI4SWhhPXVJUYsfeuIPee+R4
WGv0WUvhzWAFuo6pp6fZeuKEE0trnHl3lxkL+PWZ8KS4s1XdGTNe8+zQ9NGqya/w5d1TnFw/VWxd
HiuA7fvfeEyuRgAjA3ef0q4fk//DVC5Tsb80N87cZJIoeYXkWrBtYscoaFvQ0VzikIKaUqjO1xZg
k290YXbTnYlzDrw4TtypXjkCSYZMV4+boZZlMYgXytrONYrokW/FwqEHS6ejCzo2JHV1SACWgbbb
ptxCQkFlRu3ZGnzN/sPjqxyEzdvNDUJYrNwc/3OIbOEOpYmpSRLGicEOqxxjAcDQ2Y0ctnkdB4Zo
a6luugBZfHRCsVy8/xz8dVfU658LAs/EMhz+e951ywXiItVYAXMsFNrGRZPLGhHDNP1BX8FZrRqt
MzetbBOM6w/md7c8pElU908+4SUvvR1KD3e1SN8dnNxG9myo54AiI9gCt7+87a38jknjE1+wiwBY
LkILgvPw8svPdu91Jo5dCzsYzr0U1WoXP8fZmxxwGx9dg95bYEH+5wJn96LtVMdpVWEUQpYhvkUj
ZR6hHgzGLYbOd9MaddDrhHvrXi8SirwnKo8JaOd0aMVO4fhmZ7o7HOr9rrV27I1UiOZDkWwwPfTS
SFV9CEFDUrPikADzKQYl6m9DD2wSMAspoSpvhw/Ev3zetVDLjKuA8dLSk2pJimNINOll1tmhPHk/
gmFtmFxTy+5UL9E6BpFKdTaKNSZ9KHmcSfPRLwDGVpQBC4ili3qAsJO7/RJEGGhSTMhL1wliKoXU
M6RHOWGSh+vrx7v7FTlT5NG5Fn2NqVnJvaFXPBrR0AV2FHIzpRcthN6kyh2PLQYKpfCeMn4mrBJe
iBxNO7uy9cg3ibEzCh4uOZ2SJIAIem+p5uyIfbp6kzjyZAETtwsOzPV3KTbHeHEJ6ymceT304408
OWfmZ2wvxVwkgtqBRPwwslq3tm4uF9UiDRwEo7qUYY2vlqcu5Yc/e1JFx82yXAw38MlYWVw4lA3c
myyuPaZhL53pxgRlyLH/mq+lWR8cxNDb6fo4b1Q5XrUXqg1YJJHlKQTdwn/XAO8n2YvyFZtIZJTo
8FWOUTq1uqkMC+y45HPOYwHk7xPDAaQ6HEx/fRvoVYv3xqNRi1jvKxAgH+xFF56OOv1ejQpMu3Hz
grC46tS7+jJpn7fJlTPl3Wr7n4373LXVSPLfKokZ3bbhp5UdBTRFl2OB9DGdGEcitDuQrs/9mKz+
CjJqnhLS0w==
`protect end_protected
