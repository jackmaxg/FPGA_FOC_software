`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Kkr4ysXwwneNbLmiKAi0XkYjlAAjwEXuybA1KaS708tgCuEmIhNJCZW7ltBJQhjlZcMdC0brRQV3
YF8i8crfzg==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FXUjRWz8GADhciVAE4fmEBewwJqFOfQN5oAfwJ1bZ5rsN1OdWQXCGGKtPy7Mc+SFlHjtWcHj5yQs
zjbwPRaRwOf8oziT4rcEEC058xPKe7zIhaAKScNAXxKpdk1FHlU9A3ufiBrnevbWES5a5TpZ8IFJ
ASMQeD8u9vyLUxTDaVg=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
V2rjjnDL/QRAifL+N/57iiOGZcGGlKdVKU9OYa5BxFJG6dJ5THD1+EGWTRBuT9+vQ0iD5EwLJMaJ
TX8m6OWo8MW/Yxd5Oi3F82+kL3lbaqqzL8H/3Hgyg5pj89M5L2NNg3xqx2OIRdE4pyqBIJqWCaTy
luASMDqwiu5SksnIUe8a7It/KGcxxHt4PUt6G0EKV/5HVC78p09XTiV7C6RlXdr0B6ppd6oER8jU
TMT6x0XEQO0bckOt2KOTaO4oWiXYNjhieAu5uYRjYL5kM2EGY8LphMsq5YwNk/0BfTx6UACxGT1c
G/ZL9/l8P0I6Xe0VBF39bDrT6PfLguBD4t+FaA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lr8QL0QHkvY2RRwYKqW7sk8nUIZNq3JpVFJD+QiRjv8GEhW8JEbpsAOM2hDnwWKRpj2PKJD0GfSa
PPwnGpZQz+UpFMuwWGSbF6G7OzIRtGTbOotoY4YbypYwVuiYCIr62yY8NrOUydGs5YePi2+J6F5H
udYYL56/48/Oh+44gp82pJGyEPfDqV2mzzNoWSX2vKMz0Aos80hkkO810QTuZD2MxRhmZZz7Jb9c
vcHJqz71hj3rvxT6IWBH/asjcxdYO+xBe6aQd73sXFW/muNvho3K6ZtW66kCeSPNAd/SGxxuEjyd
MkgnqCnFg0egtGDUoreUdV5tFfj03mXi3aXdNA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LSUOXUsgLe9uZHZ5xCyiq1TXZuXPYppX9xcjIi/xFRAQrdquzzruIVQKXMb/tuh+DI01UIcN9kBL
RNXbZYPZmIEj+AHFDzTiAvPgNxtqffLUBqxwKFtBK+0we7cOGQmcEDxQoXUmsxfj7/DEnJSEJMrf
Vu8RFr6N4+5mKLE64vq66PRwSSaJw/to/cIgmBZCquMonPD4nYg4nkU8NvToZKe4/KXD9vkxijv/
Z169O6XtdlsZNGfImYmmccLmF+02slntVWh70X7Ry+gjHLplrPASmHYox+sGslF9fV85DfgroE4L
abTnnENrlJjPsRB492wOEqWIYCpB50uzHgYwsw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Eaoi25syVJoQ+vXOr1wH2LwTXhYVJsaUyCcsStHJLAbcbcriJp+KLOrOBnf1R7dNqD7u0dCiA9Qe
PZMFX/WJRjnRY+aETwvHdebn/W+F8CaDGV/NnooQgE2NK4adWfYO8vHW6qzVE4h+bOUM4StHPEwl
D+QPsAXSVUFG4GRinJ0=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
c84fsKNJgmX3tvRVOi58QcH4EGoONpILQl+W4o5A6tlc1z9zRzXB/8IcE20a6vpkdwVHWQ4aLsDa
cyKgEj7Lu8d9n+twmcyH7nklJ13EQuut0pfDjKB6GbAfagTaojObZNd6QCWtDeZESfBoE113SYEV
92imEENXVVu7mEUZqk/RbVNfUPaqdUukY/sh/zhAKhxRmZVsr8o2MDI+h9QqPXRTV7rwpK5Lwcwt
FEq+ZAbrMt8K6SmX3idZxlsaz8s6ItVzBgQsG3ugv0imubsOqDDgOC4QsQYLaYhCqYE3FkeQY142
ZiJr405Y2lI1kxs++btd4IrD/p4GNmHxRbaDjQ==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
u6onROAlsJWKsR57wU/9gLe5z1EtnbnApEmC0/11ee0/6sF2V3fDzRtngB2/N7k0PdEJT4N/0sbf
9d49iGxmWSlW76WVezmo/kA/mwnVCBzsP0EFqA/i4ndRZmVLdJuQUFFU3AycLhogmrWrGvGfgIE2
ThUodmkrBLJHSfMP3i1+Rv8GAizJ2yQpa6sUB5HXiYRG/084caijywcTzcOiC2VnV5qplEVmOXV/
pE3dUxWn/7/Z4UfgvWxhktCVbt2Gd658o+YmHl9m6Z+A3hlzZ1+juDczmCUzA3SAFlIOpEEJD8b4
jb1X/Sxh4nULtLAHqYRsTW+0GmqCxcuWv8+RBw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 133280)
`protect data_block
7N97ks9IgA/KUqUC3aPIYHDVEZmQoKW9al88kpBxOxQwM1XVGelpkh8Bw0eZhEAfppVWsaR+7nuX
AEnTcY3ESd17mdd66Z55Qx5jPp/F2VjapVP3di5Xh0N0pUD+fKCpvlXBrFL2URvHTPVaPpYLrLtG
FWxoJh6U9l9FpS2mSL/Dng+kbNc4kMWiTSOuk5ZFELI0oeapZF38WvSH0A688NZJJtJcAo1hXWZU
MCZlMQkaco1cMkHgVghnKQZIYk1YHsrS5+zQYoMXGdveczjdt9zGY9A+cbfdiaNcmkVer3DoGdWt
mJdsO8a0zGFmpmO9+5mRgAfw3o4R7tsXBWpxYSCT4kYc+RxuKkTe5oqsRVaitvAy2MnS+VnWdEt2
Ie95nmT5EcQyH+JKzh09ij8oKb/jECN7990FZbN7XZ5wNkHYALlLPf/sp3Zv6pJZf5QEFIhDFiyg
haNWZxvNh4Bm8IVTpgViVKLyuzSHhs//d9ZfuS+PnQO7sPMIcPKTHX9N64k0aZPbSKP9V3DsbCx3
RtLngEBxEHYlLfpP2o8A+TDEshsL9IqY3Ioor88I4pz58OVOOUXCGi1H0gHpEETSYSP3vPSV8eTW
c0yD7eIoxXdiluYgecLwMrgqZevzH6Qup7nASC6fJr1s4bFVLZCHK0N25Xq76ihKd8hVeoGxiVY/
xanOG9kRYpkVQXxGkAcOYF/piHBvA34L8ksTBpo7We9OrGHa/i34kFypR6BiqG8m7YpnhgASlQGR
dGjDQy+wo1EqZIRSE8F/012nLFveXEdfBGIe2FiMcU35uWWjjh1wO6E9nJbBpdxr94JMIm7WqQFc
TQd3bwPyxUePcVt5Q+4mHR8XUwvWH6fNJI5Hmh5D9ro5fowBKk1NNtDQUDq4BRzO5PD8zaA2oOz7
xrUNygrpExA6jPDVA1cmJVx/u2N+QzhHKlAGm9DMCigHGGUHVR4Nl5USWieZv+fiTnbVS56f1afI
m81fd8MGwxhssjdoEZZuUO748ALEqztzVNSytoWrEdftLW4SpRxSNv2boZ8IaNbqnvlfkuY6kIWG
viPDkq9AylfE2JXd9dGTjZjfQQMPUayA5B7Xkaapv041LE9NjTTxt+6Eu4S//MeW6mu7McJWsXhR
HIX7R5PbcdwbKOgkKCQL6NkIzCNZBs/j0LocnPPX8qoYix2dDEGn0Y21z6/7mmcJ2wimjmN/t+FX
XqCbT65HbBPR9HCo4SiFwrMi2oq1IN1G2Z2Rhq1neyg8poINFQyLfCuCyBJgJPDZunRerI0jPRkk
EBf/j2NOtbGLUcDZsnldbS+VSzzssfbLBETBtWYgIjT1vBVbkux8fjHOu5L7aGUHu4Vs2beX8vLW
Qervt3uVJl2ApUjUjky1b+DY0R63inYxFkcV2cxEb16OT8tYpRIxXRDRbqSbzuCc8S5yXF37Nnqg
KqsHPBLLs/VlniAukfFPK1TMOXo7v3+XGRrmAF4ueP3XoHe/0Y8sd3tKtrY/zJFUH1OxBF6YX2zR
zYYhP1Stf79wlQ1GPKmKR809cFYGqVpJY2/q6RWqumgWO82fYtQLmOateBT7lc9D/J1IsLyT1pbq
FOQGMtKbAwbM4bptW35OP7BKGiUXD49po5kGBwoNqWiSXM1EtMGfQdJ68MTr9yaIUw7VhKXC1UTc
5RZimQbMz6pcp5VQ/zkW5ZlQFqcogBUG9adkH66YfIFeBd1VfjQgLJi/ezPsTMgiUr+M8aWmvfJK
n5wI7ySOWs+cKMZ2mHoF+hJQ45aX/ejfeIPO4PnLTyfGJiB3M2mDrnYk5cuhrJr+UlINK4wOU6/+
jrJ/8Ob8NHYZJyot7hdH+QUJZP02X3U2051arYkLMNFwjtsnmzjqshcS77m1AReNXpyfTWOcLjPQ
HTikR1G26dVj4K0L8AGI6+5rLlFZcm/RHY5Qt1h+V/bhdi3peKihdIFWVbgddtnz6jBf3UExpz4M
qcMkSYOMCnt3+RxB68zH/6l/FmXiZQHRFcHv9UepvFJEZZ2EKkhHCDMZ7hvvM026Bl93Gvtb/2Yz
g2fPMsfaECZ8jLQXICylnOJhNqiIhW53b6vjKcZR5dL/qAmhjemHK5XwWwRvgwchejFDDv4C8vpI
X9bwZoGVTNvr6yPd6WG2q/rQ1/vYGZMDB9MhQaKnTQYaZ1kp7PK/DqkDgAw+SAVViYGP01BUzGa5
znPlcCMI6AsvHEOxELH5OzpzTUFBA+DmXBmwZlBnO8Uv0Ih1KVv3/wRFgoiNJNMjJ9Q1RDnww6Ma
r4W8DQaRWdP42uACPP/Lq6RDTa8AWH19bD67Y3yPyBVxKrAYm+Ca5JnGE6E5q8o10VCIaV+2jk6t
7DYY615PmFaFfzDoGcC5QYN6vmNeM8yTMrnB/0QtmU+9fTOt2yp/p1VhVgmHI3ay+XM/f3qBdKIc
J/ArLCicxeMkS9vKw3IOt2xuoBoyQYNHhsdabm7ExB0sTnIVkV4UqDvvjUmuIlp2EGi287bFKi+/
E8zWsb5FNe6jGnrLnoYfFkCcOTRmwBlaAlFiqD2ubIyY2Af9GYXro1r30zMFutu5Ducydfu9WIRb
hqCiiEM+MFbbhcDUutNyu95rHQlio98JUU0PW6d5NgYDx+TQpvKQpNa/cMf8LaeRI7CYN8owfrD2
8agAC8xAehdkp+kFxRqc8DDLduBMQF77GQVPl/4Jb0zgujXYp0Q92NyTSjDQR2HKzawXxxf8uoN9
nXZjWpjMqQpWHJCykbUv1cUFnPPZwcUItfjbsLYh44ohNq3E1kXwRcMImxV/pJdBgLF93aABU3kE
KfK/wGWBrr+rqY3FAkkTO+Wnq/daPMy2AESK06TGOQe5d5Z/IVKwwASC0V6Rx4xOhalIqGWuZNL1
jvDeN27Ma6UvFMQ5hZxf/8MXW396Nu5i1Wgsxg/W871kogqx2jHmrfkWatbcztrcns07a9HE6X1j
ID+7H5pH58+hYkmEh6QoVLcG2+LpJTH7qaMRJvdjpLJBaJDL8k9H4zxAzONd7kRotvTNAuZ8D6Ge
dyQldo7Dc1r8Lnqda5Y4VKuAc7j+BAXhSsQr/bhb73fw6QMpdgPVAtb2cH1bgMu/IUoa+XRfkdxX
fHdl4UAZNGU1GtXIk4NctDpXHTWx+YOZZ4czjrPFyZF5w8sQ+UonPgE6z4/WgDJ80rhbmv8xcVC0
nzXsH7vJMNDdomxTwQVCeXuStbGhPwXeXvrTY3/2sZN94annVSOpTO9gmSnLn9JgyoD86QyRhDqh
ICQIgJ4o8//GkZqs4mxlDEPFkX+TU4GgUuLScF+wnrz7glz6MypuFjMmM0z3BaJ3kf6S9/hIHsO+
0GdoGkwFUfRGemhObkfT8WBeXKO+K1fl50rfXFkecA2yPIOzdrIHLCS/kaFWhmnxaycj2QjOv5B7
6zFpeLm5BCLnjKYDFmXfxD7Zd2ua67EBkkbajxLFKjtfnoRrv/FwjHtKrSPDMUhd1L1NReTNfkWX
Az4W/G28HQfNF1Gop1G9IucPZNA4lX5Az66v9l9zclpaQN5E21VPIX8ryDxkP183psQtOrH9JB/e
l//nct1gjH9N+/w4puCt5kQBwSBWhMcuxwUGZuRKekWCJGLQ7xhg7agNZRqbdHpO6u0tA6bp2EZz
piuOJdbyuVNtaTTzQ7/lYONKRclQKU3QHlx2Le8DZIV5fq+fMyAtiVFTmJnr0Jz1eHy5FdFnr9lD
rmfvGLkWjSTMtcNqWeVbI3Yt8O/00kuht3T3wW7glvR2mZXFWLESAoJfwZoeypNbvqzrTHaLR362
5LO5sCFi3fjHu9ftDMzwaDk5jP8A5LQWU+zQq9BfRhYfgNWM37z9K2OBtb7tUwSVr5NT82jWBnSW
A7K27SvEebLZ/UUZZ+rRsbvNUoxtexxwGcwtV3KnsDCKX1SVab4JlibIS+qaQGCQy6pwloXB4r1X
KyRb5muB0gbTndqDMdXZcbPeYe8OJa7dpzeX40cHrtj2HvvNwowgJ8hmOyVhKRPF9u1uauXVh9Uz
MfZVCj5mts1eEHecR+XHhzUijPJGzWfBPLCaAPn2/Ps19NJ9eYhBbq9h+C0m5bv6WFza8jJZ8IXE
XDj66NNk+iY+OJInzkpTIuaMJBHTip9Gk2HF/utoKmWITGWVEmwwM1mqC83Kwn6GvJo/Y4r/wT2J
h0nLSyGdCiaZ2nhIgyS8kS4huEHlizNUgEUkN3h+89K+Ley+Yl0JEqik0fvt8VkutozMzueJJT3b
CkBLDQ1fyKGXv9iALgybEyMZ6NR4OYuZTyvSE7G4cVh9Lv61d8JfhxBkCm8RQjdbyH3RySMSsbEj
UlOBykTHYsiWdVpNsGswpZohsy0MLFFVrUwLIe9skgG9BOLzCuFYfUQPQIA1Me9ihOx7dvfMjM19
iEhWFh8dhilUec4vaLJtai4iC272EkeDOEhzj6jUS46EFxmF2rqLGkvP+1dDA+mqNVWn4olQaFQp
epig4oScd5TIrCA4vqQKzJ9kj7+Te6DO5Ob5m4qlNSIolYFcMNGClEKdQXFyzrNk0yPeMbD7F6d/
NM1cKzQf0jm+T11yj0Aa6BRlgQiX0L4Y6QGK0gqjrueJ5qknBV2VyIyppZF72mQXqs7bVhuSvqXu
eaKqO+6/qrtGQ0EijyPz0OINCyB1iORYmlLLVfPDN5c9W48X0XshVJcvZ3Tvg6z1cznm+aWPk4v6
KFskWJYuWdHTh/IS3Nc+2EkczBZfhE1LYo5NgEt2KxBdGO/mk5JL7Rh+K8RyoNZDBxJ+gFS1IJfB
gqqqH14nMlc7M9m3UkL/nq7SkkicLMQHAjt9DXIgADYHx5fJTiWFDhZQVg8UXWLKCNcSkNzs9u3R
4xrROEHIzQ7IRDci+clqy6SmFqxAVGIS03hRhDEGKazeE7CgZEVikMQmX7wublAlDfQqAljnOybV
epQwPiHiZmGwvozRVEe7bp8o8e12TZB3N1kfbqIfx+/sf+Vdh3hsgXNBxUvdB/b2oO6QsoEF1dge
KDTruhKvY7Evp739iFc/9RZQ8bLa4z8j97+X5pdRxVJ9c2U883lqynU0oORlxilS62EltyFbRemc
aiS0lTLHIGxjEbibIl69YZxKEXBgZfW3kdBLNj88vD84YTdAsI3omb1+P3LXxaUT9WS5k09JXTML
7UNYQ28qKKYsmUF/95e3mg4079ilXuuv3+TK/iQ3uOL993btpPMQ4Xm2UeModzoqXStix1NTDkkx
8AtrDrTu5mZIopihsBOhmT1yHSlnIYjYXgiPqWfMIvbM+edUkI5zd9QVLaTHwm9afRcajKmWqxS5
NwGBntcHZaHfd/TVvr530foBvVII1Gpx8ItwCtcrz0aaaaFBIhZ4rE57wGUYoIrGCyVTsp9Dt62F
aqzfqsIUN+ZGMmf2nz1fmcZjXhsP8nrgShzUR1qlKDPjB5FElwPmliKoQE8UUfvKeoG1aDUJpIw1
zYD8XP/ORNqAXiJTz76NTte0k99jNQ/wgFyOJ1S5oIkSwxvcnzfX64bq6RvPuplYb1vBsAV2qvMV
nAcovOmOrhXi/ip5xse4X0YITClXLhDB41UCQbYUGeW9wfP+wA5Ny2qKUisJ+tFEsazo6ksixryt
3pY20YxicsmnTcl1c8HQyKzMx9lY6wAGFNLkmxS5ao1M7rXou/Cqj5fdyy2BNA5WdngokzhqwX1e
OGHo+iomWjwuk3DVotkkl9yBC2LKl0plfw5lYYbBIcpQvPQ34Tw6lNpZTqfrIoPnYQ7J1L+s2jMV
j3h2EnoEpXLXyY3ZtSgnXGHcCrFvRQ5W5R57WToeJb74vvyyTdj9t7AYjfR8OK9gFkyCMPb5tsDn
gfbWOuM7WZUTB4eznPTuFvQiU9pyxYOkVU51mLQk9Qz4Rb6OjinOw3v4Kx8gW4+iTOstGknsnZTJ
A9uu/lh5uKvP38t1TKMPTauE1utYu7hJae4+KSqna5Wscw6VJDKx0AAKg30qK95iIo487kgzRgRh
hhdhx9KpCREAkOiwRpL1BU/A5FQrLqUgPEiIjKq6V8FD0vNOzVNu0vWnrGwUrJTbvwMwvvQM4LBq
CDRcbDE0CBGKiYC04OSgGKrSNeNsa/MKqZ7kn7fTdkr/bO9BetD1CcvskPca/PT5lfKxX4mZmxfq
L534UgVU/2Yf9RtOrnT9KDQk2GqLk/2bInFbpXNe+zYdd1bgcMvz0SKztT8Tz7fLmXF6ewecMJce
UOPCbIS6/lp/x7GQsKn+XpMfvmAMeRcYbRYEhz9fyV5au694c4baDW7xj/TY2VCpyV1um1o2h53t
bLYAYko7uIUxdGO5tBCwJg2YFb9XKf79RVC3wg8knVjluxur33kJa51kpjLelMqQjjSaxjt+uaLZ
fkvrLBScmnkGUKH8tqLcYljla9Mmi5A8G6AicXUZQu51Km/A2OvW5Vo4ENmi3C19H3G1KRBbnHRV
aBhYVmPpWWAXC+IdpvBk26nlgUf6kpLLIU3XIwgk2kTLMRtzNaux47S3Ql/HTxdgYJR25wInMQZ8
O4Iy7+tWGUGO/+tXHBeyKAir7hJMLWaZEHu68QeK5k5SHHfxZF5XG+A4qmj//rDxuLF6Fvb83Te7
GUM0zKQxmZwROzsApkN4EyEoUnoD5hRj8BRWwaCcx6F5PHlGXwkxJ2dr+Z6YoPNcE1PTLojeSnH3
euLlRoLCUa0/Ciws+xe+LjCw1vXDr2NBMhr0D9NBOv2xxS8GhQDPHXpuPo7vPljVfigIQjOH/wwl
/0QajbRpaRKltEFuYJBoHuL0e/D2GyXIJtpqfcW8RSXHrLv//F6Rx/xghsmVwgCVCtnsCSF4Nsdy
xpy4iz+sz0CNmpGE5fLrWtudWTnX7z6gckJ39dbwoQykI4yPIQO3rMZhIoZGntyfdWpkLp/VL7UK
dbG4IYN5vfmDz17X/1nrCFHVN5gRrIn+9YBcHerd+nDcjaJnw0wvNVIHZErvgrmGY7t9W2RMizoz
w/o1D0XmJboG1dBtm93/gZZAU/uKIiBgN8N12XcJD00JA2NaoHf2IjCEWKn6Fmp1PHpIX2Ip3LBP
H7xN/1/DTACynwHVSD3oxAGNGdnXzDLcXyCiMAYCaacIQiWY908NDlrvBENI5HwDOWiHyDCTgrp8
1G+uts2p3OeXQ9fLQn+PMzVSMVX6PzWypxU2KcWjxmVYDG9M/D588GGkhMMGwU4olzgGMot5b0H4
6htE4ujU9l6fqg8SZT+0AAdnADg/cYrjZ1eQKzRt6rO4V1kHLVUQrmhRgqQKjePM+gHk8o/3pYWU
twJB43q7JmodRv/Xzbt8ngNEbicIoIQyR1vH2JRHpfMK/GGWFG23hjEsWarUy8yJJ/4Gn3eLjNE1
jV8LmgEzvYTmUxOT1eoz8Yphc7EYeUIbRG/D+wCnMaRAOyMAgHvrjd8ZTj2HRNQFQH4SAYoN0X97
i7W11+dBZRNNuMoiaUrDs78xuR79e3T8xGE2he/Wy/o081hssriXsp2yS7KTGxlpkR3kTg4eC7DA
Tjc5dAajlegGLKSRj9UzBEDf4c0/7dGsD0MQSlnmUFUsEtDmHjs4RAWO1LoYVfm/GHJbuRqetxXS
MMgsU5URVvigh2/J4jc7PNlJHDd6iICo4NDUgPEEPg2aQou7TtuALRd9vhsHp+HxkOr7xEy7WAbB
7grl5/ywuZjg270vIT3pX53uZbkF+EsVd1AFn4BVEfKk0h9ve/izgVDXoKlQSIkTCFw8JdScE07w
3M6NXuATOt6Cf5/IXmU1l8SN010RUk+WJciPM3/oy0td3Tyjrko1pFDPU/F4VDNKm2asYcr3TSfp
RF4s+2yDTAdBv7Ubg0kShBpJk1RgTI2tbFV+UoxvOdRkcftPuRUdklsQIKvsfzpg5+cxHXGHgFWA
gckgfmD7efCIYmsPkyTCcCJy0QD6a+kq3GK2CsOZd9gzniqxOevf0NagQ8P61rbQE/rhlbQwjrlD
pB/Pzta6sQyFlGBGXOMkapu0VjvicewuY25ycKTLaUkeBOtUzOEwjbHzyL1c3vhx5anoGw6eqD16
iH2Vt2GkIdaF6o8J8BWZiAeJtMSsZoRU4wS/31CLmSFN3FaGNY7l2iJIIXHpaREJ4jUPe4vK9NOR
efPCqeeccgQwoTGt0W9Xmq3EDpN390uTlspW9q/F0druZFfpuHU7ZiwpIhFLdaqDfEQpn+ymbfxN
z1tVrw3pLVRFUhA4xhY5t/pejlJpidSHOFhV7YGYSvo0pUZqMOq8laKF4OP7VNEzwqQvk5fpKdPr
l+gor8cCcb4ekYjM+HtX8Y/5h611ytUE/pT4SsVmOtC4nnNrLu9OG4MTpk0sz7FPF/AQBwVtxEFM
yLbgwQN7hKJPMYSLz8GGTo0hJrwyU8tK38LTQ0IWoOe/wd2S032Bbmcu1a2eIwgoH7Kad0tg3icT
DdyJRZ/0YnoxguNQO5XMUAECXB1Kxvj3CfflmTjo/pf7vYbOiwdY6+WDQjCsPclfFoRvneeMgA/X
EokChdlud8mR0Po/ZSN2dkStK4ILdwVCiiVIRG0zAHK5mrRhG93P/CnNlPnG2rSiwddg0aPnyFc4
tbQkibfx84wiX3t9SMF6phq9HTgo37Cbi8eWbH/ooxG4hcS7wsKNMeE3N14DtEYm90TwzA1gdMAQ
ZVS4oNi8E8c+2uh0oHdgV1fMK4Wq41eNA/K1DgiZjRnExgwx0fZx+Ds53875FkrL1fOHPqm6NxZK
znQ7rydSRtdxxBNXwZX4zd05tq+EO5WlI9FB3grXFt0Y56j/lwjT4gep94z6OTIAU4+lZzYklapV
WpXEriW3ZwBlkO7GU1/Oe5Acn18L9cw5/SuuVDgHa8TBHIoeVhklnIfyWgxBdMqG5b2RvsMX/Qr2
emhFRwTAr/6DS7oEA1BV+wKRG/+Fej6NRfpO2drI2ds6Ejap1rEvFlYwxev1SOmNVeZJz0Cir2P3
OCbgCanticsWTANp3hd9h4Q1Be4q+IhK9TAeIA+7OxhEhmxmqJjfeJKhoJ2zsfZKA9+ugYnnevN6
vFLeBhdJNCrD/gHAA9DUo6EGly3GpGrNL8bI8h3jSR+kfv7PBvXWAgnbpEv/TE+OymMU6Cm0vXwF
ea4+hcUKsd0f+xLb9DcTDxKTB/JuizUoArzRI9e8nRSsxnAKlKZ3nTs1JiyDhFF3r6/xOq82jE/b
C/0ZrRuYIsc2pyJ1sZkdV2hDf/P+JaUlbVZOr+uOgMiW+KXB28XfbARJ07Mgv8vWDDBEBilXQH3S
1N5Tlc+HWsvuQcZCVl36H1mQTIwCMah85OaZiwH1SwX7IWB5npGxFZ3GuLUFF/ppTvWz0GQNYpWa
C37kpssb3nvLvaoQiRGagzCgmxUqIB4KuIIVEKLOBX1LtrWXotRDaJcj5dRroWQEoMnrn4LOWf81
93Jxxp1p5ySQ127OUJd4IQ7Yk/sXFAbyiE2ZHx/28Rg+J3lkaHgK83dsmsRs51xouE0hwX/IzdPf
9cpNWXqtxNT2Sa/Tn9OPgWonpy4Ryokw910QkJASZY1AFPFsoIAhfSmty04fmXBo1/jHHh/fd1Gk
Y3nCIFtLydnowI+mt7pJCXFzeQWbDUi1ej1LE8hPGXb6vCyjDjG/nxGzI7o7xZiQ83Ik4O7FmLvE
yO6rYGVwtRc2+24Qy9Iyl0oFqOnUick/wB+fpuflW7EK3Y+FW4Atqop/K67HmwOr9YcvKiomG9HJ
FTqV8qmWR36AGQCXwGHVpfnFHkAuO202RM0B3aCUdbvw3pp/I5aervd4Om5Dva/9ZptzPPWMoJPY
HFQzR75RV/LW4Uvl8ocUO4YFa1BEXTFh+ZDt2i3ga6JVMMTCmvE06YG3ZKnreuWntcw/B0GTkW8U
CYFFO1JNw6dC0sw9QHaqaZaXbWEihuaM/D2CK3P4RMyqozAKeBje2+M0en+olaDh3F5uSwwUUKzj
l4dY7YYvm7JoM4LB0nqbloBaJRHVQCyxZEf5BtBXF5PHiueRGmsPtto4Ygi3ap8vJbYAqTmGL1Ti
5q17pGx0S4J7F9CgHbRieutx/80ey+P5RgCgur8bEJxmXapslXlbvBA2b0ghad8CoL13zR8yDwRB
55eI3k+vivB2SL2WFUtQUkqRqdB+O9owwrs6doOB83Lo7k36zjaCdcsdkOaJ98C6KnV4y9xcX6D8
P3HiGIfbM8MHvFIamHy/ilUXzrb8Il/XZH5N52GuFUgePPxTZgiV5H+frZ0/l7RcpKssIz6meuSa
2GmzWXNwaZoeaNmrmkui0/QTUHQtEymeQUvGp6EqWrrQToPbmb/GIGLe5p3dg9Ov4/W9XABa3Jvo
y48NLoqJf8mD3OfxiZtSkrg9ZRwjQToWrS4hFM4XSYkvNczU8/dDcQWUzMU+3khoRuS2BQcIQ3j9
ZjD6P0iTl35fA//OxIougRK93mi8G+OkT4PtD+DM0X8oPE+Tw9Qq+Ot2huiTS7TD1WEXQDPZXVQn
1PxT+SoVyvHox5xZr2VpKy8a0ZcV4J0FYo2Pd6U/1+uOUqB1USfn5uC6mUiCEluV65kFMzOgxbJo
7fBAHufjkEws3+pDCyd6TJjGVck0NvkyNbPoeqiMl+za6CVV9QGE0pizsMKqD9QJM2stczg3+6J7
cBNgbGHcHWYlbf5A4jbb+pVlFiBoRSJ/Mu2oUCyBZYmifFGmjsxMnC6K7daWFIfQ8MnfZ/miW58X
qudUDWdpeLQh7188cil3Jv8EfGc8Dr8M96syEQUyu7YtNKy9cySEptnRwRLIKnMcR+/JyRFc9mKs
BkCbf75sodqoUAqSZdV+5QEqp+0ndhE8iCSNv/cB/KG6o2Ymfl5bnR00VzyLxafYYndjOVAQH1uJ
pz/X7AW1Wb3g6XhcDouRomt2vkAqMNkZTTT2yn2s1cE6H3CQoX7EgXiaCe1+27YKiESoZ5O43Xwl
thOdtCRVy8InJbZdV41/cuDAKP3UglMHi8yKVBeflXQsSYDji+5F9/AMW7K51u2o0QofLeknYGAw
XA/cOLewNUifMEuSIa3/I+nOgItTaaq/+q5M5W/7FkNyLAZ/hl5C6shwEKkjUC0pN6IzvzZgN2IX
fSiFRGRoacuUbQocAIt5RHZfY09U2uUZ/yv/JImXFQM1zmIoePf4XxPvCiAoSnPOy8AWP/q2cKkv
VWPBKNdn3Q9EGYIOdUrLjZ3u6ediKApZhWzFJLBpdSO+Uq2NYgfnkquufJmg/Rt1LClSnZGzsTXt
jTcoryALpwu4kIuMpKx5QMnrGqj2RckH/o7eP1QhoBaiWUursME+C+JfR/9B6oWofkdj4sVdUXfY
5SZHodrHuRj7RhBlS3/GtOaOMEJgy9ZRs+EGdD1qaVU8MplJpZ4mG3rHeiTjfwOK4UOX084sz/PA
ygbA4e0bKLOm0jE4F3fq5gtPD8EDBcDKtX7tZFE7D6q5qvZhstxxOBj099ehEzpveC100O9ddymB
LQ1NdEzBfyqxpVLYv2027tPS7m1cI9wyOmYZqmedqKgvPgpIvRKtF27RHk3BPInOzuVfEJr493hu
epcQuLrXkpyov7WnrzgB0fxlJ5xHNlZVdrJDpyGmOxM+i9Jn0Skg6HwTe4RdDMK/eTcKVWqaQPk3
272/y48tlFgSVCAVBYxKPLGGxnY1L+LhEQ/29WfHaSaT4eQiS2k4nFLxKBxjBKNMCzp/gTiv8i6e
qCgahucgVEew5AoK3zH6CjOYKYwLV2R/VEYHBSvxk88oF64dNoca5NnJjOH8hIvxSYWdC60LYTio
C3Oq20GpEC7ANtdIdorbCqwuwPUJco1cIJohqCkkBv7zEY3yNT/nwffVdVuir7XDSCo1l34kd6xQ
H3i6DSLrJ/fwEUjevES8ZbfdWXYgYAK9/ParlxVmB3aQJwoLM+XTvCjK+Dg81Xo/S8elTFNLbpE9
DqpEmoSStfCvUsscnEn9zlzY9adjkIzjUR3mRkVSqjHELspx2TTxbZMrYUFsTpxN1S7SvoTPs8/B
pGDQt5niPC+hbPzivi3zoQWdg6jkgOpgEEjJg7FD05C34ylh6xtiHnD+w5YySS4+GdiT4YXEDMtG
hDFKB6ledSASan9fi6/XhSNGsbOUWSyz1/roDT53ma9VJG737BseN62h7bwBwXQgMokdq1L/AWqW
+gs0TfdtByjyltpFkURx6d8DQ/pMx4yyxYsHg3uTHKl+W42fvaINDsrPBlpJ49gx7bOtr3+VBqYT
2bqUz+ouEUkvUSnTGc/r6dlIFo2vgc8uvQDwkqt6huFQJufCHPD0s3/u4vvFLcmh1Vw9X/OxlON7
ax7xeA+e4UH8v/mydnbbCkjaRLpUd7E0K9EXBqMu5EbqsYOovO5HR6cMNwrYIRnqSUm9plsYyVvs
8GE59eTFs4NEGYyUTqHkvU0j8C4eAclfUqNaDbCovzPgUUeCBGPFgjCTtP7HbqpmKQT2MyEclXPR
DPrOv/pnkIsmn5OyqOM41SE2xrjXz3NWHX9FXlnete9yeiGN90k6HBP70cRHThQbVlJj98pibT9i
p89Q2OyMLQigYbfXbuNqnsAEXKPXNeP5Stzdb+Q2GHb2BU3F2ttmAiBixuEMbEzDyxRHvSb29BhN
0AdJeJyH8CCUnsx916zcbLl1PYZThC2Ty0aqw5d7Ad4jVcM0py8dc6FLum6rT02XYVvYf/Tftet5
G2phz6AfNf+NxsI0+LDwKYQT7JmNk9QYmbHjv52lxyXK6i6MnykOaXi0+GdCoTpq4daA0XqEVFZq
YRBmAKerDHgPXrlOSGwv2nIgexOss7exIacmnqIaOxdleiQvEsIa7ZVQ+p9RqeWwqMjvufkwafRi
bWuehfYaN8xxDXjJLQ0TQgmljfWS7epBj5LwzzBFgkoi8PT2J0ChjhCNpprpsgro+B5jYs2xp4t+
1+jWZEHJZcDINSvZ2JGp47ey/H9cDWuNs9vuQdmoBnZXt1DXPp2/9l6W/4vn42NXY71cOQIzmO4D
ghcnu86CrnAmie0mVZbhEBBd81wOx7tOFprX944HpVZpIT7l0MdEWxrpT86m3HwglMClLQm+46Pn
DJF1XpNEkgcBo33L//YrkhdlFAkpGeyMBMTtXJfdcmhl5/+7b4R7Niwf4Hu270PGrXg5mlFfLutP
5VIEzRYI6IXrvVP9itdBjX+wmMstp+snYrmsG93noeryIBMFvSfJbIsnS4u2cJtlQWop+ELi/bHU
EwTBbctGxXtL3CqUB4wiX+Erdi/eNp3WN9nK5+e8puTOuLuE/WrWfqMR/KA1wZgouZGH3+Trjf/Y
4zZaHJbycWcVlrNsups2d+Ocj+QULgHraEsyirOOIlKu9bApGIkRZjVIHSYz5oC4LT8eWVr8P2sP
41v8/AzBAK8PRCvQXJC1hQFocGDhYJQE0+quKId1BNgvzOtNZ+IjiIY7SUhSvjpbKlnekRL5xghN
txnmdEfG8qKK6DsTL5AICwHksbnue5gv7m2jXb1cTHTQze+sPSGVHwy79VLd/tO/muVYamsYPdIe
m2oNrQxjTX3h0nashTr+Inec7aAkgfHjBQ6Sa5t0xK9xohYL98Z2WUmvQbshQNhiIPgC5S+QdxqG
fWTnf72LefeqPkNwuX0SVO4iR1imF2IrwNxy7XMenVvqjYTscT4lzlzFH40KDfLPkjLzoX20gA9J
/betsoI3Pm9D6BxKhlFwd5GB8yD4DpI4FeXDkLeJELSZqkVKrhRQRzE957UttyCK6U22f9SOXgIX
zP5520CQb0N3ho0bwGd1c4yDRtxT0HRYw2Po2YBdMJ6ZGiLLuxR5usb6UtId4pnDJdHFOBcnnYNJ
vY8khy3Hmos/HCCQf7r+pCQFBPmvjX7uc11pjeA2oK5gik9WphogebZ+CxeB2cyVf78kkL/uPRUT
ZA+S95qvEXMbiZnpATVkXWgHaPQBhZSw2wlaR2xwk/DrStPFCnSmMHiS/ESvfxr6KN+aw2mZIss/
NMu1mmdsbmc5amxHTrhzeP4pP5tV5Gn58WW9A2SYglTD+8Tb635rc9dfhNGfqcivRhw/hX4lCE5g
ET7uiBXIuezj5WtkDAb2JzxnUM4EVAZW+uOuLUSETpMcEeC4nXAwv/YvUPPA0lmHAaL+62HwNFoE
BoEdRhvT//pTBsVQqz7WuPzpIzDPG/ldLIFpyTtDWMnrccdIxTPjh7vaon1TgVDivX1TSNrBaQxn
RFzDsb1hcQe5NgwvWnjF+U6zsTVs7qDkURQKkkdxkkrcig1KkyWfK3jFiG29iou3LfJJsaAU6SFV
a7AxXNIwrACa7wGCNW4+0BEtvAli4owoq1sqBTZ8nTBwBTk8+n9+sJVLuAbnFE/Y7134aYnwYs9A
ng8yWwoRgGWRS0zcbfVdH63SuURNWvvuIyWUu4knv8hvBICEitPSxs6Ux73YkB9lWPz1NHd4slJi
6hG2cJDIw9der+/3R0dGOMlvhtwvIrN9bSOd7NaEUd9V9m/6bRMgBmWsnZtIZvZNjH3gN5uasfkF
4iwwdBVXMMqvmz4VY1V3/JAM0XE5HuGiPhs5uLAhTZtk0jatJ7rGkbXq3QZsxbVK3SeXG+sq1xOG
UeaPGEcy2cj3Yj7/xhaPs8qcP+XqavIonP58wW8vf94xF4a+fmgoSGF/nTWYCFuvI9LpmzmpqyvE
1PUktlcl5xyvdIt59jtMPzNFtvJ22WcYIemar6l3yF+HCtex9ZMZtOky5XtQ78AMpfkUyKoHQ4Ow
2/iUrDyxjN6PVIfy6F83U4NunwQ1tgIN7HXnvJPiI0jFGj9OmPRZOcJW9qqaKoGAIUg8oEB8xTJh
F2fdIdkvh61SE73LuzIn5hzXo5tqa9fxoi22Xx8JEyPVS7rwHGDahQQa2HhjJCjg0Ponpqxi0s2d
dk9aSquN3BkB1R940fuY2/Sj4YAsxL/d9IZZPVeLSM/it3YDi2Qg+uUwxXiT2eNQyjhf4erapCNL
+8D1l2bCKU67as202be/y2rLjJWkVD83QDDopqpqHpHelKrefh4+ns358xp2tHWkb8MhotbbSnrz
NHdEzS9aPPTmTmIFPK1EXQ0JL/V5JozbYmoBgKx98kgQ6GlsXrk19MkB8gPgHaA0dr43HsDNwFyB
i+urqtF7PIUapg2s1GtI7Ons+LiOhHN6NHJD7dAu3ALTAYO8DQvHSQ20vaaoEVC2SdqSp9mYcunE
Xyc2iTsW6N3zb2dOqeJjORiu7s9Q6m8WqmZeMXEZ0B0ib0T134HMZUe0rsOq51Ll6ml977VceWaY
O12jVzizpyctwOW3XH5YxlhAe4AJVMrmcq8wTk8ykh72rYND5HUkok3U7QdQJTP/58nZ0VfmFf+/
yVsvfHCeEFm8W3KIM5J24g1JeWK1u9wDkSC+hHv/PGEwyFjA/x2ZVCwSYMZVwWVDvde38M6DdUDd
dIew/jLJu45UsDJsAcY7D7dU6AKCEpMl7aR2mC3y7f8O0CW08/SiiWu2M5ucmt95Mh710iuLZVwu
bbcQAA+ceU6E3R7nAipXeCFBVbJgBWS6jJTAt/tYII/ggn9aCJq06MGHqoUuOM1dXdaIl6vho8Nx
pVbZPGLfj9X8pu3fIIqjiGAZA5a1YxY+nPMIJ75PKxtkMnlXFhaXD7/p38+hpSe3vdfecnAlX5xl
WdR/8gvpU+EhiOc3ysj4XhhY5MgVObiZrcZdpZ6NsLnfnWOToeI6yuQpIiedVauF/E/2sTXvW1Qq
Md2lTxu5+tkiHzGYYj4IeUT83oRTapnEuiPDI907aNg/RlT8n07gr1ihIxwYb2zW1a5f1b/LDu2Q
062oYfcZxXYZwstuB19jyLLXrAJ2fUlc+yVFR+uy1QBEmEdl6YkRel7x+dOvIwHnBe1AC5gkbFOJ
XmT7Trd50e03dV/3cOTvV9mLZtGf6Rg5XLXIzZUQptxBmwVly0bQVKt/FJg0jOpTL2ngVIrLVp4A
mqLtwXT6ONQjMxcb3E/1jCNSLvM4Fa41dBrz4G2zumh3gfl7+TKSOAIHtGc7VAZxS5+yEqYl+Yt9
VB04uXKMRpSztkTIBKZ3ijTn42pSgS+B4Efc5kj+VlayK04kliM0b3z8AaXv42eayIK9+w9YN2iH
RassVPu0EVrj2Tq+7cs2rwtVwt7s00Ihtcj+vGBChOgz7yi9YMjRwrFd+K+ugHCGQV02NC0Uq5Fx
fOepYKgZSbhVG2h7LzIw5RKcyUnOtCHjaPOyNGgYkZuOfr1iOAq33ZU+eyhzSdbDgY7bZeds2YAb
+nKRlMkwxSJA3mNOfqxos39df5p2Ex11GpCcTG2GvVTlRH81I0FqkcgyEw1whUWExhYkl8aruob6
RxIGCbNeZCoPgNoCNleqm/VyLBjxrmMj1Y3u5lU7G0+Rk751MG/+iXhee8h6t0XVcsquPCrGUKLG
9NCarD2MPRPoyAPbX0KV0yVDdhDEokD9nas3WZRVsfQdu7Eg9ITyELi2LEfNcRgYrPqahMqZw4KH
80fkXj5i8VZ5EcWCmofO5jn3ZcaoDqiVVYI3JqxovnIFLMT0E9e2eczHCiagW8VhkMJ7BfvsQllx
BtpS+UAD8rSdTsSgc0TUYoEitfHQ4kbLT1tw4NnFLvlSHkqnkWPntMfInbkOGiEp0tR1Z9SnOpY6
oqiYOHAfrJhXaEl6skpKNyMQ1OD4cubDmpSMTxkkngqASqtc5wUWq+xV6tC6Z1ynA/ZpBoyFERF7
/a0xeO5NUzpfG6TJLvrGdgy+CjX+j4IqglZ4aDCIGGyLWRG2uGUbrRgmYimp5lzlzCRCPVwQ5FhM
i6zEi8Y+Jf/cDAWye34qaLlzIm9YsUzXVEjz4jderH6B4ZNh8lf/C18wSHw62GiH2RUfyRxp4jyT
SW9/eHde+WeUekRqx99Xo42i5M3bWUHg8M/noNxVFWyrjQzV6hz20QMJeHlsJ3yo4wrGLV+8D5pU
Yk4wjLpsJ86z37Vwa8ydyqCT6o7mO3Xqaqrc0l9Kdd0/DY4cGEr7ocENMKm1qdymDaBx76HzTTlr
CCoS8MevFUtJ+6z6Tsyq9G9Ab0bX1GX46h6t3Ynq/qZ3ZOiYj8k/zXweqm4YU76wyoMQnj7AF0Pm
e8tMFJbLtBJMgT2urYWIZkf7c7avCgaxpkEXPLlJSRnr5Z4Ug3XySDGplEiCE6QMFw0JE4V/MBg/
z8sy6ZQhDxv+lLq8hyNFOh5nP+8iRpAQydRCHo0qhnaExPuYfzeoqupH4hjN1m3XrnJaDPLeNNzI
kB93dWFiYYRcstAlvaE+RYVJFQXg+ixq3BP03xzjJeK4r4DScSOe8i3KsbJdTzD+dgfrc5XfEqdB
Gxqbzs8+wGYKm7U6k6LYroEvq8oLiuLn72Dyd2y4afS9be4WygWGxe5RUuGObDQ0yD8byqi+eJe3
yOlwoJDIltAK6JU3RYinlYpPGj/rFodraWYr1EC81mR2CtcFEa7L35lrUvFTlhPel2BeV5K0vSLO
fA+q6r/RN52UeCgcThqInChaaUW88Eri2yYn6apvmBTIxufPBVjG3lIK0qwwDv0NrR0LOLAQa9Qi
EJVnY6mJfhqztCfjWbGXk8/kbgA52LV323BQ/UehLaqElX1rAsyeJMQycaoBCwggxTxgm87f0GyQ
CEugRvw3cJgrmZrCaoRUvYoJqA7GLh1A/JWybyg/L4aGS7iPOULVCW1GIwr7twTl30RwsFGpAq2G
rL4xVgS01XjMSxFAk2CNpqZZUyETWdT75DpCWWt+CZDES45e4ym8Col9X7cipg9L9ff8dMS1mzWj
0IvSUgpdboo4FUX6qEz/Bd3XiHExfB+5myov9Jf/t5FrBNuBmj8Ld9cYyu1Y96TMEHSqCceb10Gb
nFyIrWjkF06+xl339ySm2GsaY5TzDTyV6eVO3UnNmv55HjNCK/yOz+cM4ODixUt8smNPJUK4i9bK
SnhM9tWvWbH6qgqoQyg0L9barudQe4WkoZTBl6K+tflxe7LGsoDFU/Re0Ztvusjks5H9WQCexkUU
LePpe9ofzORP3r4hAJLOms1zopCp+GLSJxUQ3OpyLqumQos6FK7m3Yz5HqYWnyvQLAu1naYv4RVG
gHOUfRIoIPvr76E7ssvIlCHdJrU+SZsZNcuCmJ2R8m8LsZkfg5rA5xGXWBb4raIL08d7g/O6WRCw
Y4lCWhPqM33LMu0STQ3jXxxkfovROvRb3pYvZWpZuqDT6r+2vY5cqEt+DgjiRVyTzan10mV7U3Pf
UO1ltYT60aqE0tJnaFb8YGctuMxb5vnbhfRDMsZnfS/XhdpqIXHoCLunY62xA9nXBzxqQm0G6R7n
fLghUVWDPPjWbz/byCnx0UBeoTUmwFOy9+XNAdGN514/UqN9DcdzCaO3BbhfTXkzrC608zqc56nx
6NSEjhIZvsEaAox4kElZORbO/LRdiIIX5HpHDh3MQuCZzA8Du7/BBihnP42MXMIYecyyGfM3Vqok
B43N9ZGvl4lTU6UG0Io+MhVcJO2d5FKB0llZS9ucHZXI46X2DAXWX8tl0Eb47ISU/GEFHdDEwE4p
k//iiTOHiHZyyPLyfGBDF0C0UxkPh6x560826Q6GrGpJaCsT0/qNe8UJfOBZ50jPHfh620teTr2G
5OvqpXjQTJuYACIMiva4L8MMk+aKlM7TBivqrB5a+5Lr9ApvNPJJIfXyW1hwWgOHT4iUe2q8sBkF
R6OGdrV5/N8ju8qpvjSDY6MzY8hn9CBCAZepdOENVDckBtGQF/jh4gS/uJQ5H2i0QR1vMo7+UL6F
2ww58V1Jj2/FbASELdsPEkG4YZmkY1AdtfVTOEFDt3W/Sf8BkrUiq9QSXmWHtopLBnWserDPn0xv
EXodS8hQZau+1+KML4Nj7DoDtjgetDwulCsymDqKpqeahCstOfu4qgbPJ1Zalc0++8xgL2r2F2WF
0iovD336+nGhmXrSrFafa+8DODETbSQvmynLsN/9VGpiLfcasXZxAi5jmDdGna69FTeIZ+jwjSaD
Pf8qqlBVfULZ4oyI3yDRAKDJqEn+X8lxLpOQbi4PZdum+yTAo2+AAUQ5HbW+4yxUQH2NsaIAS8gz
hi5FVQjRoytLx5jL/539NsArmYE4zIi2FB4NOTJ2f2Gz37+AhdUs/j8NNk7gob5DB0LVpeSFM+Zk
p3rjdH7AuYkxxy7ePx405qXvdwR+mDECa+ativMGOC/TXnBM7wuAgmv/KSOrhOZa3GAsqaDFkXWB
mXqjOLfdfu2xNZrDAy9qi9v/jO8PgIkYpzuSeQI/aWZ3dolOhXV7+ACXJyq/oWzCd176aTntxipH
a5/UDbg+fEKoRKVCIf1Xu4Uzcczt+IY/f8NEvGVNPX0vPcJR5gdrkQQHh9G4mXOjfyjgCdCCHo38
Low5XLiE3LlgIIheaVIP4UVY9HVRPf9lPp5OPvH/+YjWFvzU/ZywOK/Zt2vd5asIgdypvK9SlFf/
dzhbMQWXiPFHgdHtUWnIewfo4G1N1W+dIQh5YnGUkqTwoJ+xSGbOMebX3j+D3VC0lcULvxoTMfuD
gSEULH5kn10YNMNRvLj5HT4ptLyNRF/9ZMgrp7I36VNlMuN+x/RIn8yy5Py0343yuJyKOO92ArKG
4njGyQz8bpavTzg8Piw0DSrhYhpEfnHnZCYczf1m9IL2e1hsxY9VwA5tmUSXLxgvHrYoOuWG2jZB
pCULtNz5fDIm14Ef0pA0oqNdcaIOIulBUgJY5pVkN2/RZUajeBt4DxgMg8UhH4RJIgCjUZ2jzcg2
jO3sY/bCfC3TfSDfFLsjAvPgTZGWLFP/10v+qMiAW+1WOGGdHb8S+zXsHLiv19pHyW9PBQJo3Xz1
eLPQEzWHAiYf4Ws5R/8rhP583YHvdj6ZLk2vqitA5hMxnugCXGV/L+FiMEAJbNEPC6yrJWbRTLI6
B8ZTK0ONstGswVahCy0wWr8UiYSjOH5T0hqoplRd3hEZW19X68bmI59HYD3bk8aAUUL0opBzwQDp
pT8LW1KmY65cPzskxfOJ45b5odDsGYlZbGMdYWLT6DOlAUap/ggdZigLbd54Z2ORHzhkTn+JlnDN
lBxC3ZcvkwohC7URZ1n2li1ism/nkG7UpRrPTMcYEOjnZ2X3QdNCUl5VanO6jJeb09avxj+HaJ//
whwjTloQ3H3cfDbQCpY1xLmqJ2pcWZ5pRHb5xzGF9m4jU1Tziu0BY/85rEFhJxlLG7aSbkZ7VAxe
TjxFEl5rE5i5jiAMnE8Z2ciJ+phHt54a9eWt3oTrVIdrJTexZn88VD7x0Xhb/0SoDXrKwKixtjj9
SIvUoSoWYjokuLmxP2GrUmpi7Xec6HZF/fd7ytC3WkJNvzFfVjeXSp+6n8phVwZy6pqAnE+hzrJJ
trkFCEvCAS8kB9UkTZApPK9gaVyMuqBsNSHEOXYcr95QQJu7kIXMIPYg5mPrtiQf1C9B/J9m8uXz
Ryqb6BA9NnMVMfslo+u8OOLFBMTKaCeAsamCIdPrl4xM871GhaJ8lpHDeAi2wJU6XLbibYe729D4
hJzQ8Kk8x15IUD3JFnSoq/R7rFfIcuSrfg0ygmn86zbo6mD83x/gNlr79xlHmrzOoNPdViwl3FYD
563RvKimOTHyXgiCf4pobqQgbbcVAT1+hySaeonvs32XGP9iedqAk6LNmFLZx175fD4vrgmuSWRO
t1A4nn4uzilGTSnXLiI0B6uFVGS2qUGoBxLgGB1y3r8Xq5t+VLPyGmkLhUAqAkABWki6c42diF7Y
e1jjObXvsyNv8jDGkO0fENb9hngtOaaMpRGDfZAwO8R0jaLsJezi7URdQNg+5v8+O/6Q+P00Tloj
bitbAJp0e8joKsNAqfjG0ZM24dgOFo1REk7wGc6oIrNNKw+zY29RpEiiZHntzkaCPDG1IF3mtvSn
mG5Rs4FwkyibIhvc/hqT2SRjZP8j9za/A/1U+iip0xHn6JVes2sFC1BH/o8i4WmGxGY32fJgXlPg
YwaEu1+wRFRGPWEVS6NS3MSZiGzhEa89xdCCtjc2rIjV+kSwwmQ0qx3ic+8aGbO1hlWQsviiRH+x
IHkLRZotD+gtxUsSrcqKfOcfIpUKAAlm9sIfxkbhJTT6ZLsvJODAuhoxcgC2TgCZX8BjCbiFXFi0
dUlBz14CKO/cl4LBzEG6bHxzcU/GUA/mONrSMKPM4UICvUNPf3ICVJVBGVcD77Gh0HER/fCa2G04
FVVsbAbHIn1dgMe1TdptN452whslyDlq6Oixle9OyOfeEXHgx0G9yLCu9k2fdDXwCz7VjWiy8fGu
W0RRDcoJqYtjktptZBjZIu7ZeHOHw8BzFeVhochMPujsjqKAA2ipHgWeVioQB2HSTpbs0EJlolqB
1PugrfOLCT56lS2qWtNuKSoU/AsL3XaWvycDLD8E20afiEU5JgbtoKDEubR5QGAiJKDjdaYFYA8W
R6mFCoNM17VXXqeE0OuTqcZVt2ej6KZGpEdB+lm7cLnlcXgndadsyyHsvOwUiulCjl0LEfZOhMH6
nlxi5mU6Frpg2hpkGzCDhxyvU+qxLEtKPzQW+eLOVFDp8qBgHSvfNodol1yN6uDlVhFrqb2kNxyM
7n/iTSLA9Bqm5Ss3l2QkRhFJMcOfnmmcz00iNoc8bhgR7QKSwgT3ZorjGciBTSeq6WbSiU85OfP7
ZjpwvDvmIIjPEPl00Ha0PfJa7veWETdqeVUp5+hRYPdbcCJi7jh9Eo5oklD/JZheTUlY4IM5PjIW
Sw78xzqw0Ga5ML+xNjnSA/zJtrjBI/fqOlI0Mgac6Jj15rEBtKj10rB4+VjGbdYlQ5gTbxjfTVEH
D2ft2wOpJXG94IDt4G6PHL+iKzjQBwg9hp8delGYt7+5SC2B2RHBfiq4DcX+Munoz4jw8T7Y8VKZ
Yrds3nJkzKsq04uHUsKbpsls0L+ktIcHs7Otx2q9mPX1uUjQf7gw9RlV79RGo9SejnAGvOO7/gCh
3lDvFJqBXH9Lv0ADcDVbJz4bIpWPsPMnWrOrmB6np4SwF34QTC/x9d3BaUVjPhdCfkcWLlTh87fd
zXSI7xuFJv1VoywD8otRPc2Qx5f4WH3AlWvaFriezzMnopKOSyA2RexawZHzzL1Wrs51GcAsNS4g
aYbYuy30fO1iMjBSHcLtHPIxKl1zPnJixTMv9OBmkLXB7Z2KaTZVE+OmMomcx0dZnY4aRQLnpKH0
CN6zc1Iy/nh7PaAPxQZ2Am2qEmouNV1lxSbLIC230Ub2sXvmOjRUFP1xbHWZv9VypODpYciG5LUK
O9OWhfaLEqRo6iJF+qS9CeWsGXF4IMD96KkI9HT6C8A/xyl0TRkCG6V81qYzo+5BCWS3A3uOrpW8
4gHGSWAQqYkPVLejWWkjrTvq8HqqYB7LoB0mb6uf81wQV8oLasQFid5kjMNYBWyHRCwRixTsN2Ij
lJDupsWwzlFrqk0SH+zJUOhz1RLCfsWvHRHqddCy2KuTxO+l2DJb6QUlaCAWaMpK/0hWCUSPt3Wo
eDiJmZBiyvBPRtbukkxHe/K6kl9BO0smkvQlNSI1Oyy6t72rTeZNeBDlccNFMciwQXV0SD6P1bKq
Bst3w9s4ctYTsJ3wn53kijfalLHBGrU43xN65IFIfbb5gmti2RdYKIMskWItjodNdRLL/rqwDTU1
tq20WZv1VpcFT0fHBRz/AdsDp0P1OSX02I4ZzE3VPi6VEvS4MvOrGtKiSNy8rAG82l0WJmRocJmD
JsQjwgrYow/bi6Z+eQTcmYPkrx+9haI4TuUGp/n8oJoij/Qo0zlIaczEm4alVO6zFxuBQD67tBOI
zZlyWIl83gL2r2K14N+AtG49QHq5iIDa8zeV2t53pMyjVaOkfOM6bB+tQfBrfmDgLffsVpD3mnXg
smDyGNRAkYTiXCh3wpHhjfCagaHfiohKEksaYbzrBz8Pg3rjyttydQlAbty59U481s9/Ec65P7mG
yzXy+zuup5uHCIzcuv1ZreikCnRk4RSq/Tig7vEpIsHDjRuZxB+g/JM2ZnNmm2Fcf2wu7Y9FanQi
tsm8g72pdsDae6msZmzMBtXAPPZwYAKWs0DvuX3NRz/fgHu66AzYFyw2rqLvcZj4HRO6O9F4Gxy6
aiICK4MCsOgovgd03h9FcIXJshcLSsTwVVK18JEkNWmOe+k89b4fYpX6pN2SS9VRtITjabWulykP
MkLwqB3sdzi49UvTnrwyhkUj0bXk0IhfT48LWsdUmWQ1xUTYwT6hUooLfmGiJotxjhR1Jy3PFOct
hgdGqB4ze0JHkRGBlcQVWh+aTU832SnaI9WM9igdPrUUWx0fZnRdN5Vi30BMPMp9D+tlT6LWlZSd
XNbbFqz8w8//m5YmkC1hn0MPPZKe6Pcx7EFXi06RU6cUtHVgVLzeswDynHWkP61UMq5LoArEyUzC
DCop0FRTF56/kHIUEOIfdDFd2uUb/xNw7SPTyWlKtKVBCQmA+JBGShQlP3J0F/iFNauLrZjIVw8i
8c7XwINjBKdDridkqc2P5eEDvqu/kKescVZRSYvsN6SHAR5C06+6eRypN4XKX2s3zqKwGb29rEKj
sFVjejQZ4ePGUejHGcmEBFeICzDUJ5J1vSCiv/SMCNNdRA1llzM8QFAI3lityTOzrQ9GGXAJ+uEE
MZt33xjHtmoQN/VdcWh8MuxmAP84M/B6MEp66kLRR3N+EIJrgZr8oRO4PPDnWzjlpQqyeT5TaVQr
i48EjWwPKlkA8xbFfxB6folW9gsGzMOebkj8ducKlpYu6ggnLkL/CDJxwt0Qyn7uV4uDISzimqxK
/GiYFS+UDRvl7SN7BfcD6JT1W+b06gRCSLTWyEC6qOA/Jf04S5/zB2pEWV17WS1E17nSpLpkyhtG
XDBkmvlnV/CqxvcfV77Et6A6KRdFw5NIUnK5X47n08NjMHcJu7wUWJ/qhnHJjqOmm2JDo4wZ8Xmq
mt3kex3B5HktCZFFVDrcE/rsT7gxsOCqoJDZzblrBiFZL/o3mP+EswNBaYfEwRsQRxmvv0Q5Nh/w
EVyeHSzYb25p3svuCYkGZdUPMFEPBP090OydhrWQA0sCORgRuZZKxvQjYG5R5bINxce73pGWFOIT
AfWoKRGMUb1YO/zFhhhturf/Ew4qBsH9j+CV7KhtpX/yUkRMeWzS3Dxw99hf2yEGq27kLpbwfoeU
OV+Q4x4bUNjFTcyqEwiBJcmz7xh90QY5o/I8uqaaxJYi8HeYJqaLfADjwb5B0+Kn8SLhbye88GtH
i2Q269jmJdX8KwjQYqVwWurMl8wXHAgzWthe7pEMBG1YQQp6gTynTmDyAw8zDQngoA5VBK1SWqV9
gEYBP5YrCKRoXNxYZNl4sIVdW/axYMoaRw9gJH0dXJ/W3tdaxkHVS7p4S8IZQAyuiww+YHJTPtwI
pOUF7P4R1dCpO7zq1QmwbAdZL2eaDwc9Lni1STCE/NVTzUkT0DH2u2Z3Jb1P8NF9qblgiptAeDzs
qp1/iAuLWTEQB82guoD1FLzaZ39Kp+83u/+kf9yXL3xjwzpBsFg+WRzb9DtN6fDcvmM+EdmRjX43
A8ZamSiaXCb9CbGH/n6y+wDsRi8uc4CcsfQX0/HTY66pdRBQzJtYI6U8fzvnGMSpRDHxZ7d5vviz
YYoGNzgIQ9t/ks/PpAZQLhG2Nzm1LJtOlFog0S0en1WUy74709QzGdSNyjnvlL159AB+om1HSABM
yzXbzjJMq/tS+RybNkxMTWcgW/3MDzxfMrujgFQ0UleO08+HuI3zQk0KPSuL7z+4LLoZIueSybNb
T4TKT9qFJXIpvrBihuN1xs8lSyfy6uj2I8PxG9KdxKcO3FpdHJdeJS5ET1OFF2Tzej6DpzeWAGBm
nYjC7bcrofRcMCf7gP8NGYveqMaKynA68Da82hnBET9qDyW1SSlh0gdB/ZRaEqSU1iuN519JQLHS
C67E2V3dQYLkYm3nIk4OMgGAgavTff1hpelmjsjgTGqhhgi2J/sKdg8FC2JS5K/kcwQglnXcN1k4
mgjrrfjdZHLeXRGSZ9ffH775YqE4GPkaL2vOTF1hw4mRKHJCLD77Dpwejg8F6Mg82ppNq6xBfy3D
6FKLtrKVF4+wW9TEzkL4ze5ZfssiR7zyBn/Dc/ROhDB/DzRNg7D/udongl0exXCOQeMRFUc0RM36
mAsW6IQtjNPC+7Ffu4JMqJDRavfbt0WW4nyNTspCdM+2Z2QAVsiW4EUdzTTQS9pVgi8Zu9BMG+CL
t8BE8jeG2JDYZX9hAJyBaAdyKqrS2Yq5eV2a1og+H7+mSxBOsMe9BYJ31nUspQ8oSn6/poc53b7C
MO6zvMNTTv1cRYO+90sKT8N2XuVds0U0ydblWcyXwIhJyV9DOsLfvXVrFRChBOwpR+HQtjquT7eQ
sZNtCfc3jHJdgCxxYA8lLYE+Q8pdPYihNSDucV1Go0gK4EyeLG1pUNd0amzvbRvNkTxEZk+PvR7e
Vjkgi3TOG6hben8kIgabjaC8jlrdMtHSBuEZGURtk0c2XPEac7++2JubefBme22cgQxgEZzNHnwe
DvK04wNKzpxgE6l7d5ujQIJhCGc71P+hJHUcSKVegj6m1wDyC3ItrQfFuKPeG6whCwCKAcyOBdfY
Eo56Dh7/I6USsk2a3Ujk+qysDW47dUMX8C0EW6Q0eRZqdHoe+ddODq9F1OyhKnDKAqhhokcbBEG5
6v6gq1bPvCV0zMa04tcYOOvaQCq1+f7y5YfoyP9gJc3rIT3xKgt3SSdfLZWLJy1z+hHTIRUmmcuM
1NPc/t0Jc84gLlt5dWXSVagymg4Hr975mwwW4QLPFDpnkD1EcTe8DaTEut05etBMz9SEzXL3WINA
+sv9gt+7uE8i9mx9Y/j8sdLhaDhHBBSHOa40P4UeMEhZybhLNA5JLqNJqbVzNCWOFjoFx0YeLYlV
EI7M2+MHz4Gmfk7IJ2ODQYJ5/ztY+aqoWCVv9nidpfuZBUisJNDic071APZLKfynNWjFGcS2Fqg2
fCrLRimRzilEh1JuONft4Q+SxwjcqR95FJJN8amPQgO/SbiWqz4RtXvlMnuqwCSoGDukvvT0iSRd
LxwFXcoq8In0a5gLQY91u5OlchMCrnPmJ0s6532Zg60D+98lFrckHuKrgeDwT7ltaSPKSsy1t3ZH
VSLlFcGv2n0cJKPbtbrAu3zQykkTkG1/ATNS5XexxvRnF0pZx7wPikuJLSICKTOGWdYreXefDmYW
GPXPVJyYXbzdh9RU4qLegs/gslSwd6WhDTxD0BLPH8FA1nJh7KB1uIYc1jY7be2DLtw+rah8mPNj
JYGt8qVaC/gjBq4nm0hJJJa1vVeoSIN9xh3v9KXUzMBvBJWX6cH5gUNr3NxWpskdXT6EE+P3cYqf
G5dpTFjCHmqLxbSfNu9UdGd06mlkevkFhxBzQ0Ng3OS5QhFBCTFtFgH27hcrt2hSKZ8GJPLCzXat
Bz8FIiClerp2qtCnTVGyJ8D2bL6dTYn+wzxsLLrsHxrpadsKjs8ZtHKct4QPN5HBvxNhKTwIqIVv
NxI2uoq2FlGOPi7M2Pehd0OTLZsU616yGzbmJ3saw+UOWMm1WDZ0Al4xcSKYN2dds8w+S3X/IynT
UnbrCSagG6WyVBmpZxyxvGl/wj7xppCvfmqMbZL1hAh+w3tkPiFyPthpkbf6Aw/we7bQl7xNTiSd
fC7Tl1mTzGMCmFpo3IkajGeK8JLPEoJ/9zHZhnZiGvyuOSl9MXez6jBXsRkPcSleDnJS0hObtOHK
+VYMd+T3B/iwmmgjOiC/uR4XjNMN8XHCsxUnei9Wt3hq1hIaY4rbA/kmDXeItDx5E69W7h1tlz73
/EkzjvppMo/gy9vR73JnYKq3G9HnY6xcIUL8CSxLNVyZkeBmgpuXBjhStVoANvtUoqPeLtmNmLfD
vVhzwjarY9egd0ymRgSbMH19VzUT6OgEj0NKoU/k7/ASo18ydub4vhmMIQpOvzpXchVciVPKJyDT
7eyE7Fkd2i733ah9uG27ocqtHTejR5GiH3gbYLTSHw5T3e9f9Kess7K3YMGd2BJZ/aGcrBMecvfo
KpZA/rd2fIo0ODcdhbGzM7GkGShYwE5stMFdgJXsOj4u6tgR0mk7dvqK9MfiLl389JTRFP0BMbxW
L289RtU+08thdTHWSqZDcJlpmUYMEosIDVEwWGs7VO/YbiL+6g8Fgxf2qUmnNpo4Oz0Uk1bD0sWG
lcvqc6jMOb7yT1Y8KtzmkgpNXoMFd9XAoDyLV7GnL2S2Y+pMrKzafuIt/OEWEaGES/mCkvDNqo82
fOb+p/gHrslnhlolkI1GUqau6o8YChn7Tq78rqx2sJxz1xiNN9vpk/JVllRlAjoEMkcMKirqlBQu
moV8RFoyPM1RmDeHVEIxukngPROzzI4OshFMS5raWmIMLX4rdy08NyL7j3KYLxclCs/FQZF9m2Ec
idVqJhwhunaQx1exdO6ZQDa5RzqthJQnbHwhkOHphJC7/Q3emit0qEdc58+9cgI/b3NT4wXZTbPS
sCkNCXsGJxgvRh+ttOU+4fI4PJpb6AEc99hDNWkode552vcZAE44+IwXC9zvmxLa2ocU4RQGiSh6
agUK0cmmLjfAM1h++Ty7H4uMRvxjnvsRXpyWb927ncpgZbmrNRMtP1T54nVM1G1kPlwWZFKZnzbq
yPFzhdKWOg8n9LvggExrpGwU3xaAJ9YzKkdoqX00Ss5arIA9zQ8EZwHTC5ZdbeHKdiV3ucrjxCa5
q345DKTa648u2bGwFLlxWlgS9iNWsR3GL08OScRRlCOwHbr2jCCtaEFtJS4mX1kA0P9pPNZk/xUl
0H3kuwp/DiG2NfWRKkc+wIjVNx98fBd2L+hqljcWFjsWjQFylx+IsysjUCsiqTi8LA+JFKwiZPN6
d76fc84sDI4Cq8+kuqZX7ZcGXKnVuRE+6yC+aUxThmtz+0cZAaL60MCU8CeCPUwcVon8GzRcXar2
2RVxVn6FZkT8Zu+95WxD5wo0xuerSYzR0yvOsNjjekH9aik/T8Gc5xX9DcP6IOEoS8QGLeJi9/dH
CidZEq+E0Oj6vkyrxxiJp9Yc9k8Te0Q8RZhEUQyWRxEA1WgIhIrrageUIeGyxSxxGhvr5+/QR/cK
1Qbisul49LwXDYO1xSTWw5p9LirLp1kRClLpCqIE4Jdd5fLsmhmDdRdOouISC2/w1ua7eqsJq9LK
Iz1uykTkKsghUgXAPkktmQ9BLFacBlEsx6Ax5fo1eHA4HS7l+VwbdXbss6kyGpF9szCjqpVY5NoZ
WzVwd51wF9GSOT2favpxm2VuWXOa0nhGyccj2EbZgxVHDeMJQRfUGkh7gbzV+fNotHdh5EYBow1s
jveHlzUatCyC1wCkgGMV5Qxly/uYkdTwffBUP9Yvrt30rJXmt8aTPQbNS/273qd3RwJfSPWowADE
DH4BMteQZzjOhI1h4qFpm4T0DM7j/QU4YRtr+7eWbF8pgeM3eSafuA6YZjydF4KO+XJbe5HvfsXd
hNZ1+ImtD0VmaJmni7GP48AlADgATxEjxFO2qE0wyNBZZiciR5GVmk2gOREqlcnsPa5bT+kYxUGc
txNSUCfgehhf6/72cMucgCTJN+4TihvUeMYpu7uLpmPkGddQuK95OeR8ZMOoEsOFkucojsa61FNC
OeCMbqC14NX1D+YthB2I7KIJel7QUNvVXOw2ugxAQxyOekmZUuE6oknjh7EnN0HqlkDsgHVGTyue
dR9oqfaHryOlEmoh+IgK6XYTCrZnKtaTxSrO364Rwf5VYQ9xBXLRc4QcKPq3V3Vyl3IStARgHeXj
6VQPFnfY+xmPL+vjYctoUpeAP97TVyaOA21S0NLqM3nvw3oHT4DyUmbnMhN9y18tidxBA73feEYO
B9bzsYl8j18OCc1fI+EoxMNTXZrhgWFKwrTXzZgmg1GApbeDnapw3KczWIUxHashX/V+cJJBTids
UXX59tJxmuqa409a96VZ3AjDMYmhYiwQEz4xUYBfBXYgDNDzzVP2huB6IZsdqlE/gkcRSh55xfsQ
LHBrScaT23e+P0miY/JUCC88I0qn/qiXiH/2eVJSiaFMPikWS4MctBAClgsAIoxalPMWOPEWXi+W
CC+BtdmlLIeeDpiN1PlAtonTaM3bXXKrwDSnWc2rsupM1KkfX15iathXf9mGfXx1E6JYGYQD6AxY
JlVnstBmpCt/ZV26uQFLYZWHKtC8DmSSqygIa9SZxLyQcndqwoT0i+l6o3TURcp6LPGNMjlPy/f5
QJLFaijs8BJ1V/pAkvEX/wtZ+zNnVOCM/alM+NQ4qbWge5PXVXzXWYWndJsU9bpRQOIXqJX7W82R
VlE3TBDWiVLQKxXMz5ETEjkOwTH2Yl4dC0U72QsSLuioLv5QdVk/554l9NVwnrKwBbI+gHhWe6sD
5YJbh+gvVfaBPPlxqUlpoKUM2xYgRvwYEJbBP0BWWhDA8ekkPP2UyH94zdr4eY9xXb+zU76HDgR1
Q5sysGk9/VIlK2NTaEb7yYQJHy7uafrmWSPuaTbgb9+lQPnahFGqs6ikvEzbPF0STerAPm95H/rJ
+eeNbIpyBFk20og1FLJb9FsuY3rU6ohmvR2JGiWeHfx2vOPuRtXLSXy64ADFHMZhoeJTpftk9hY8
6gzLq/NebR4tgr0e1AQkR4xvoGnwyK+gyPQbL25TLOdP2iegnhTrMvs8INrLWYlAkcuHwwGEN1/n
fIO3UWna/d/XLX/bpZnEVOp5Xla7NYHIjpCaAJ+tPhI5y+I0LFprfDODju7bvYdylJ653bOg+tm8
GZ66GN324U9YmX6ryJxGWWjJsyaKTyLvXbTyWChKuiRrsGAe9JupwQemwrdADzdI2RmoMS3pYVMX
aI5fK3F71EorxulpSqOwiO363dQglTiz7zdFhkZ8oxkW2rdDLAV7tFm8p0nj7sERibGSbdVN5T4e
+FtiPmAewfxwYfJVa8sTdDJ2E5C4wCCZShb+Rq7eH4d4D6h5ABzBdUAOCeRbmEXslZSyp4PqC/G3
qf8g7cG3M7pSvL6e1UNExIjkHvpfw3HHy4qFKbOpGYzoAlSHsR4Q0ch1iJkbL4jwTc/qeJG2vol4
EGLm7E/eBHjtafA1r74l+CCautWod38o8e6FEdSOV8Qf7LhBSjKexvB+7xB9L34EOroBT7LPi1rj
yOWjkAgzXmEqHizRFjuqFZC+xbqiKKUSMfyxyr+kfpcAdrqY2b17YbMNtmZREVmIYZrZha7dAs6g
Lv3pzqefCHlbWIc9nYSfwBmV8TWzqZzuSsEuNyrj95pH34zhprva2AHKD5Jt4ZcsqDKhMOaefhNB
br6IMvdpQ2hIEizfHWq0VLJr32oc0Ny8VI8VdtHL/moBwVN6/LXUygdlwLiZ6f+qWUJJN+Rj574S
fiOqBsLFLSBZrDesK5pIVhY5u/2iD+7IggF0n6KWdAIT4n7K6sSLkXi//JjUh5wIW+Bkwem6VDmO
YaalZ8KVflgzpqTG329sGt23tPrNbfklpc0EUkfLHugONyggMPcuSwsHQhpqTbPLGxbN5fxn5V7/
8WzFAxXiES33OWbQNxftAH6tf0SYtfftOsfsSV+WzD9Lmql1GMcMYTR+sVrfSU4ET070aZ30jm42
PtI8gEeE548rF/uzzkoJhfFR8MuyV70P6jCzRCpDwoHm3hiLMAlEasOH4xRGplhNKS1SUKzeWXH4
PEnKNti50nzZEp2NTcqscziAW5YlDVagZ0FcifyOhv5PmPhsdavXflsj3+D++dz88KcrAfUrm2kB
oXgnaRyHxH5JEbeJzOsHbUBaweafYckEFUAEGfQlEqhlIox8+QC45i6cU9VUqqFvt2VBTdRQeCdT
VQ/YHX6llh5N8OR4dqUD9GMJwIZuE85w3chwQRDZA/0IIwNDqunkYjRMY5GjspTtGBQPA1AkGHpH
RxHhtvBnyKlgbEWUqoPJUCS73DGLsmJGcDzkFcdJzOempYZoOIEMhpv2Idc0nWpU/KSBzz63Zzjb
tgB5xM3FC8fijKzLM82qw2pZTGHgJC5w4XbH5p+KPrvP0eQ2q6L9kOrsdiNqz4oHS1eZoJt+4/EO
AZ3xPLzhMuyabUDIbq+HKfR+mocREU94q1+qpsGXu0JQO41/FhDGLy/dO4Kdd3TKkqE+mDzvaaOT
X6CwD83ujYkCNVsH30zX1K4zVmma1D6r5v/1fDS852m5Ggvx/wHQulySw1QgYoktHS/BJGUAMWtv
moEgeBtiuy56e9pMOIocTrf/qw2rblsaSSMhb/q3FZ/t+ZbLeB2Si3IqzhMEOh64PnjdKrardbv5
87Lttb2JY0BWDYR+siWfr7QBK7+RM3JGuu7I03IwQjoKKD6ToRzq0AjTyLEoL8bTsNkvjM7ltv+3
lOcqKSoXQ45TmVFqOaztXL2Fei8R1rB2gW3EGDiQjS6HlucmgAzZo6LP2IhSvAOOqgp0I8+TNv8M
syZerXYSU/0jMwNA+ecY2Am7z2beXSR5fnUDgLJQYgHER7ji/pgF2eFhxB4VAwjfZ25W4WaQ3UcD
sBjyZkp2dgGnXC+KN/S/NKMnu5wcTrLIpCP2wQ7RXUQ4lWcnuM3GqJZ3fIGV+lnIjWh6xdypc9pY
MIf1hW08Zk+A/dQuLcVoIabeMmbbm+Qqpogrmm2zajMBzIb7sm3XxYV/lCkL/i6pyPHprEy9Wxbg
uVxJXklGC9xsFe+dy+7eFN5bnmZs0li1XyV8E9mS/jYr6/kClJvpU98R1x3yWz3nAkqoJ9TuODQq
EpWF7LrerNKEIoGb7abuxZNediG0aiXKVpLDjEFcOBDhCphrwBrSSDistjRqsA8I1CSMtzMzDMtG
dnF0vZxtdvMKNCda/XfUzEtYjpKvvPNbNIxeb8Si5hOCmAJwyo53Wc+4auRItONsRD+ZNPy9RZjk
RU3t4d0Q0bBrz4R+wOAlu8kujOpxrDGpoRm4mPhmQvGEQkz1G40YKkgjjdszYjd90QVH5FoRAuoX
7OJTTeKjc48fx+f9VXHDUlQZkXvGKlOl/aXzCFH3HJiXfeNtIOUdK8FQoS/eh0U+1TXZf17LXou/
JDBl23JfhBeJFY9gnwGJAJHlxQ29ZuILtOOqnz3TdAWynKS3wx4+8tWt5IR1R6hlLvtYT4+tcZ7f
Wpm+drVcmLq0Hgysmt2nz9Rtky2kouVnY94oAUu3iXDmZcliIGa+ZOJRWT6JvaeT5uRbkH9aVhDV
uLUQtAC/sCj/3tllDiQomRXIpOtT+1n5rqqDNcWyulHrEmkPSaQwztbHyrrFGCaZi4ZQhWh1Whih
OnBlzXBGG1SARREP5jq5fwU4i4MeUwkhYT5KDZ1bhmvzLJxFc5L9JnpW1Ua/A/tpIm0468wSWh+k
hy6xBMCAcpOATLmxqRkx/L7w/oC4Hy6x4X2N6akAt0Y0QP7st7biacvuVLyFRn9jGMVOHfmVoGOD
KfQVjTpM1enVx2VsOZHCcKUviR68ihE4g4DpiHh2C9OL+yVj7yItdWIwBwI7aZ9V+5rmrkdq2vXO
KJDXhANLp9VcmywNUJxvAUl9SiyS0FIGthUBGvhaq07/A4oqgyKQ5um1MM1MRGVvb5ePziF/r+hi
20sZu51tiVHMbQ3GowObIy0eBPPXXwt0nwuQZB/+saKL8I60169YneVpfMbJ/K/IsQxVp52QvB0y
615PdcaKzRHloNfAcaDTUU58bYI7z//N+I5eG5f7ZqJ1y4oy0nLtND0eKK9utA3Krzhmf/1PCJgs
RiNif8mVKNSBAGbcF/WK5kPYm3nzQMYIJaqWZOFhtY/UMpgFNnF4btQCKtjXHaBYcB3HgYCK52s7
uD3eOjxG0k11Fmx7rxrBxN1FMk8tuhbb91PiuxqHByz9R50QV8kfHZ3MwMY9liN0pKCmIeviIAfS
ntG4d/kIQzGAKLVNCua34C4y4mUp5aQ6tleoW7KqiZQW7OJBh5a5O5+OBenClqlIPyfL/Lp5Mtg/
50l/H3J6JuOPiYcawoBXeExd6z/mW4rs9Wczmr7D2WcZAbZ+n53vfAm1cgUpt1CdCDRKenOUPjAO
dejYDfjqJp1FCSj8k3JERS2GrIrceqOF5w7pG8jxE5q7C5UpUzukJPBAWDj8LbiTmO7xoCiUpQYu
GXnNq1ck/fzjVr9xIo0rYSEY5a9qOp5+HBqJDJOHPM+2LdX0AqxD499Salnb8njp7zkKileYTSKO
0wwEpyhNAuSxDwGKw37Ligu7c8lgG90u+4TNIbqorZ1QwivOjj8n/SdZqTS5b/Y2fqRDknNB/EtA
Vc33u4VWvvBKabjUCAO6qs8m3snd0VoBaDpqBNBq5J9EnNo4jYwLRjKXqcrXbxWQzafPzsKW9Sze
+xJiGAICDOgbpEShQzgws/sBem8fZaomaItk6yKCFmc3B+MnGI5A9tT/yuR41bY/tNgFwu3Tg4vQ
eD7Fy3n3MGmxLRIAl3CZKZd39+dxI2u1r9DfSbag+cxTTwRZt4lHAwkM9GGvI0lYUyHyA+1Ucq3/
wkV9dtmXqEvet6OcpwAQF8EV0nrqlrGPb2B4oVp1JTi9yrbRDj62hCSKBExCN+vnz8xtFMCCNjEy
Wkj+E+7ekXiBZiPTGsQYfDNC8jrrkCFcLQ20Xq5dlVY6eQsCc6lPrrhbkxBSAbbULJhRwVHPSeyI
2MNyu/UypsZKsP5jFlCl2jPLdp1JMLFakMWZCCRCe3foGFvpWlN3zN2jendxbewwAwosL3FFd5qQ
7abn8if8/Zk0H9N93HrNnyHVDcxXAeE5JEBVM6p6T7y5fnQJIHNQMPiwz3yWZ/XnknNEA3N9DHaS
wRr1lEP4WIfIK83m9cLvo7cAJYw7NTBaNzBcJlI+lxjHMdv0YCuh49XFe16dHA0Yw3HtsBU4O37F
dYdjjHnlm4KwcXlLQgg/FS2bkLWDuJasyxF2Q6/2HXtOXEjT9hTIThElInNcTKXe1b5BJZnNKDuo
sxgFqa2qzxyvWc5GDLtRf9aRHFXNNSbiaExZY7Oub67FeeFYdhB1RGHpBVIy/+qDAXFZyfAcFuH4
4xIhlTUborQGYy3l8Pezw+X7OQueUJa5ohYSpW5ezdK+y+/GCDMwhdTeGMTg5EyyLiEu3L0JILd/
YsoMwX5GOUX+JzZqF9QKQZNFNHyain8yzuX6LUpcoLGt/2GvzqWbKT3BpyWktIr8oIhLAmKHkR6x
z94onp1eG7uRr1z180JOuPrsutlrfkOOETWtoQqfV3SH9E1mGL+Kn8ybnGSz/DZjnlDO+Qt/QuyB
4t7cAJeW6KACIV1Ouh/bbYgY9QWP24P6jb29diwVJjDNv/nX7Y/Ig+/Y/emLheWGlBqlf++P+wSy
R81DCC5NlZfnfwbboN1WwCMx9UbSeZXec7u1Bpa2sGJhKEfdbOsI6pISBXONdhGf+Z1YmXSh55PY
SOIYgx2LQg1vwseDJqv/cKAZA77tM9z4uHneSmyhCSSZt8YNOx4SfOIpJl+1qFcBqs5QFI7pmfb1
yt1Nz7S1p5a1SrldlA6I7vJHuUtskVkFCbAYG2JOZgFIzVjl53jpvsGMCdP4oi5/FjniS81/AKrW
rHanJPk7kkXuf2hSwL1RVsXahCdrv5DyKAW66ori4qSdpSdOSYtDwLNNID9/fsmm/HnunZQUskir
W8sktpUXgHqJ/Ty9IPzQL1CC+RNRmR+hTazVP33mvYXZAxA/qEerBoW+8tbKzkSaYBUs47pdkzeo
jUbBD5yKRJ4+O+uc1HRr79n+7+BABf0GSUUGSC0vyxiyXv7hayFl+J43bg7c3oi44gjHGl5NrqUg
lGUqNcYjw3/NEm+skNqNewinOJNy28qK/Fss422+WsIqxSxzj+m1OaUtz63KQ0qKVMZCwRjSPsr9
ygikMXrlqqR8KcNhx0Adtt2yDQqbzI4a9NJN7qZ03m/FMTHf6UNKWJ1w6blGa49wSkS3m+iwPtnO
cO060b00x3k1dYLNAfS5R8GisKKxk4j+mdTlkKC5pzYWWVE79oowPuus27EwtvEE+/hniE3z10og
2LShAYQQ1gNOm8G8tS8nNxbgs7yr/7h48omVtGQohydhD/I2POnVdg0RY/qq1gHSD9ksZg13l3Cg
LON2MI+AH6eJJvG+Tpct9hOh1EiAFeeGvUsj0/HAI9ySOCZ0is/U+uBz16ueK2xneO8nBRHepSef
IU8Ilbrf+vLMjgWVs9LvW6LIlCH6zRcxT9Z8pagUvFANK+lDarVK+FsOv01HjsA4KvMXwuGbNBIr
pNyM4/PxhOIyJ1Tgt01mpfkim7MJvR5lODwRYDYPwPzo3yZv1kKWvl+s/CVyoybzwl04/rdWZ3tC
R64UC8E2DWrjm3JndOqltTEk9cE5wC/Vdw6w3GmnN4fd/+LzksMrwGgBSY6pKw+osOucgtPjldVt
Mycok2LhkbWpqUx/ioPqGF677Uq+nrAglgZtvevddaBdLY+dqKJMdZ7B/Oj9TSTpkGTkcJExV3ju
FJPF6qDQ0M+FGD0+H6A+cMnPZOPxhsYhVA0fKzPXZp2LOOzcn+BnqoxZiRP5G8Si15rnMSN0/KS6
SqvhqQopb+Cq0EXCjwef7K1e1pHRBjN6dQQ1tFsR+NmqZDyEPsJvNOwnRfw2m86uc+10A0YMO1XA
loAMWH2DxfTvYbkNnH9ZvECI7Fq9CtxuKgWSMjew8EslLpVfZ3gj+7IuuT1s3BrxRxtMTDcYR/QF
6gmbzfvU5cH8OcMGZRkI+QWT8lctk8scMNKonbiRJAAxfHU8gTxNXo7EP2byfysi6uI02w+NdSj2
z9xOr9IZK3UWoBFBFkh70/haI83egDSHNfCKe/QM+Yfs73AcSery+7vl49RqoepSdpgaEftM45xt
Wp1ab7CRvM4RLwkV+7d2nR/lWuAIelayOjxBk4f2WHceNZ1eHTJ14EVEOaw4/Z8OsImZp2Qq5f/6
qovYTZl1KeXsV55tZwoANj3e7dDUsU6/Nx+l1Cz2fH+hNjW78eZRJ9zqvDqT5NDLzkuwAxJARfn3
V5Cf2iohn8We1YBwpju8ndEfCLeCmwRKojRrlJWqM2BlNcKb3YqibINs/0ZXRV0MG45Y3Wj8Gwyr
IAqCJcJ2j0DxZ5IO6YTwyF++OF8glaAoyFfYbaqm2x3Z9FIJa+tEjEr2pTsAYczPybL7di+rfXS0
T3XZvhYZO6+BDor+2nYFPFwHoMQcqEhq3IPEdh6aLlBtJ/2Mq+0K6d+xHJSEAOa9C7AKGeqH34Oq
jKoD6G4xYBLrhbm1yvpvQ9qjUUdibcujj7j2EdxAWMdA3/tHTQc587Yz/vJj899BdPJB5Yjj/Z07
Qx5AphJdIFf7/ni4MWHeozvfQO4kH/AoSG25KXAWIqBUWcEZ7LetdMLgnONhEkmJbzKyOcsNV+OX
Xt9Jzgh+ZZM8izgeqglmPb+AOCteN0BMBAtWzdGtLjkMP28PPxqjBcvnqVm0/UbkjAHdaNbLBjtj
LMZML2UWGQ4YwE3e2ps9laqG91+p9HNwiXS6NWSog+9jucex+Jq2Vtp56D7itB4ceFsIjGh/eDfu
f3RjbMX1GrrMYpjO6DL11SWzTG2HRPwVyyhx5uwPYdXhyBoywg7IXy53U5zZrbFIUSPN9SA1Jdx6
C47hpvhawuAGZ43wF4QeadWVJWUg8Pg8zSleufpFILr/sxuzX4JuvNjr9Da036EJeCBLro5ANocG
KeYbzcUjCyUUq7IBXLiKt2gPHokvq8MrBZkeIgM2H2cfNm17FFpE749zT+lF6/6fhogG+wXwY7Ck
uW8tM+Obw+yNkwNEqltDVEG4SxbT/Mr4yj20jvOjKvpdlSapgnftgYp14lfh+uYWGkqmvAqoeP6s
nIYGGJa+72Tzy1+Sd4b12Y5bHNqS50NNSrTapLmsu7OSpA0AEuCEEcLawc+APTOMRFV4lh8Sb/qK
W5tuQ5LPvQ5dYeEllNfJXvI6NzC3mVAzrq3uGnX1PHNZBpGk/JvPjv9+CL3gS6iru3zNAgj6jK7v
m7Wvv5HHyTFbQQvj6anmEPkZ84ikmtnpAhcskBMrq00OHka+OsOamYdmZ/FWzYTUC7IgRdpq8gWo
Ru5GEj+IJaVMVKxp5c/SNmNTsewquUW3NN0S6VwFGFdaC1GzfmUZha/tJHMvTNcGn8EIrTWVPdth
BMmBQfeZOtVtkUcP1kjEGXkER1iS4xAYSVCTBFYj/S5v5xkW7soC6wajfv9Hwlj2Yc3oSZDtXXSp
+a9icW4JeGceSz122vRP/wXVEShPY6/JJEOo4C57u2fANjRgxQf6cJXpthfvhj0qX/1lU9GEGgV+
x7aqmP1EvtWAy45TVG2Mq2xCqFkG3xZIJQSXHQUxaLwHG2L0GJOvlVlaY6kaQ2qk/Koo4uwhtVPc
zbbDkVs4Z0ObIuM4quc9PFhDfsnTQZgwRedQkiShkHJVSMYFpyjn8DfUSVguDIe756CwgrU+5Oj1
xq1g49zKnDwt4C1pkEZsIL6907Kd4ohi3yeXNzOCh9Xgj5IJLAE7mFTkpI2EyPhv7zYdpeyAbOX7
Mwhp2npQ/uBNl3C3JGUqtr3BejAmSTuPQYL3mTfzFIbV/T1VT//nEbW6uQwSCEvLSER0XN/8Af+f
UY++VVHeKbcgXexgBnBrweTPk/Ud4itWB4JJuoxB9y24prOG4Amgs7hTEqPVge0gcADmFlxgRBPC
BQ6m4nfwCr5WoPdnPaUxYp+KO2Ln9pxUXLnhAccewMO3VZj2Bty15JPJyAkLkDbOXg6/1pznrlxF
Gc0QDR2bl0ha0la5pccxKLE97MxtZIdRKLx9uxsNgsF0vcJJydrHQzCJTeKV0BhLsT3GipRk5eYG
/m+YsAZq3+SE4Hevk5tXsUrKcWtVE9OmfJkkrauDn0EZUKnPpoc7Sr6ixsmEeN+fhgeh0mhuopVw
nAkgDdL7E7LzLuWbIThMiQ5mdlczzFexG8izVCV973ghZWB9SZRQ0/ZWvuhJ7cdZA2+nE9ox2svO
aKjVxPc486E8zjxcP/XHef2On1+wapAdBPLAExDyWgqgzlYHB+hZUB02EE5HNpbVN04qyaYXjb9H
1CVnpGc1iABLIO/pQcRhfSjF814WtoDUoL3cJzPzbUPhYK0oXV8fhKXz5gzuAyDGXdm7ZUscWRS3
bXVRY8eoNUQW6VyQQxXCsSCgSb4zSYx8DeHnIC4jX6oTARZcujDmnW3ukhzyxMgRVIFpukH1p5sI
byQXv1k3cAhnpWZanWnR26U6f/FAi2C3mvUK4ujxgAjE96w8UlH8AthEbAgbvzqqNUYp7ATrih3p
U0Tg7/M4cO5YZWGyfykueOGooLh0QIXiQHO/JTMpvkb5Ee4QwaTPDp+H3+zhJOaMDbZetHDY9Y3p
0Yh7szIP3Wd9PDilzAL5UMynaR+EE90uqOpcPArCsxkva5vtL9syOxR3M/BSAnR5Ej6tuw90DzFq
/S/TFWnUw5Lzumlp+iAn7HpUKp0OvYKq7OS4dw9+1+u0xqOgTthRSwvNZGyRPY1jjqN6iNXAKzl/
7RuAjIhQInIhiZLmDsq32yo2Dp9dWGuAs8potDXptC/mh6YM/rGx/maAuZu1E7bKXBthROqQXL4E
wPR51JShwWNdp4GHOXMMfOmghpXxuIpPV9K5/GAwzMpp07ZNIT0h/Jd21Y30hL1Psp+XD14BWEfF
ErYXOxLo/kyFSANvdd4UhGjqqkl3leDrypWZnB4ZB77BCMAktaEuTvgGdeYfsBuSdZ1VuPYdyY1R
6zsK3+wjKOWZS3daMvWqClitPOgtsp3QBPEyApID7Xt9b1ZJm7kpxQ2dJoMGqH4ZX3HpYRuVEIcx
tDLjygk+yp6aVo8QJYgucNNyCKMshJhT/Wbszk5jT1jcPEGqg0JM9f2mIgzgocSyOaODbXw8HKCf
59WmDFTKHOPnmMlS0MAQVBVoJyYnDrGJzo9CIoYRteJBqfxa+gvanwqxT8zKh0PJNC1nADVQpUPY
lHGEyIG4Cgg+VcGfhSiyCKhiBy6Z5rCd/AHzhvuI5VEKad6G/Uw1NiiQ4iA0wL5SCc5XaTxcdBaJ
3kDsR2BIgtRRDLnDFdoQGmjlSm3kCbU7+9eo3f1Qe4t6QRjpYxemDbFmI6abrSBjB/EfYOK5UZYc
OF6DO8UBOdJJSAsU04zpawsHwHpY3NnTu6Eaxgq/vlTVXSwelN+Jm4ETFdzDJbb6VKc7ECzj0Y2o
pKHToDwy3aCG+qHOdgUJsxrfkfR/vyu30sBwztGtiLalHXKhd6FfV2Lgj+3/4JmWbVbTZP+hQJN8
/6tgZftGxhvdy7y8k/iB6ZgqYt8HJaTBDjfjdcfF/k5jHRCLQrrPL38y+rnamoLpNJBA0opjvEqx
Trt/pC4zfQQlVkM95KuTPjg35Vb3tfBOw98IeopLIYQHZBZveWO3Y8wyXdEiopuB+/pw3ye1wyCU
3neUkV9RvBeHNJB4fGWra6p32J5RdksQO5/PJMtGPKSUctBwArLzQj7j8QM/hT0ebFkkO32leMmr
8DVvplKydAlItcFevJ3WoyRkJ+eQKuN3p1QtP9m08woRVMGf5Xz+ICXdc0DdxdYZYBhk0fe5e8N5
I9ISTPjL5EpB37O4jWxOgk/yannbEL208rg7HcToPJ5TWFXCHIbU7A/4SzJLQ2IJQktwlMR5zd5U
r2ZAUPltSHDftMOTILm8bqexNiS8TC0bOn0+631TMaURWwi7oYz8WSUIq+9PO5yQAj6UOXWOQJTM
uWcJsRc+GZ/uUM3oQ8D6Gf86uMB4bbAjFuQoqE0J6C4CYzYUVvl5oI3l2RXK2T2Z+JS73aiE43Xy
rXX7IggcKEMz5jMHt21QutfgQwUg2RaX8On2fXrlNnDyIR/vfN/+qNTkNRxrcw2VnMWIOiANuYO/
IJZHFoXK+1OCEIHTXD59PBnR6yYiXfzmf1plxq6Hkd0ulY8fvIQQXwscnutL5eiQAVHQpRxOGyv3
MMnfRGeW+3tadXQ3jTmJ94iZEbS2Ej2EEzfwsQtp+1UYMcu3pvbWuXhCc0JbTwn7hI+fuYd7ijjY
8S5RYjPZrHCcfk/Jk8wSy4svY1c6pvLeNYqXzMJega6FOx/WcrhrUlX3Fu4oD8AYEIgM94QVzgyy
K9EUmxZ0R9JZNgfHuQ7GXrESfO5NRfRKX2Cc/iBTgc8LHybrgp6ZlXVAraStsqkbDQku7EfxYoJT
Nc8t3GiiKzA40KKXPeNCTi68BbuZNjU5eIj9uK2VKx50F6S91euWvA0iAKXeEwrCL+t1VyxMzXBS
IG/+M0khBONNEvbqxZ7nIlX4xX4dtoL1dw6Xw6rOds3A9L5qyB+NR8WEHcH5N5QKvMuPBV7LeYMN
35WcybkQN4aE0vdMVPeBEznjgw4Ca4LbPP2rrXWq9xSJQeNeWgRbWTiByCiunfW9D1x8M9rqe//N
kI/pnl28pGyMVggQehkwdakNII3nQb3IDDSdL322qKqJoFU17CB3/xViBVWNAc0hKFP5CfQpZT8Y
XADSV/VsVrmltI3BPhxrwixp7Kak/+BYrk8YhbZVknjmC3x1Xfqu26CrZlgtKdcFPiNaZYPGY0zy
0hH104ARAByYj03h1kvlDMwrIhDOfi2FoxAQ9HlJBQSimpVhHP5jccV83CDdyH+ufEhcIQbtS0la
HplLON1+JZjINsZqS+JxUhjjXEt8w1Ev1pgYJUuXvZVZGmXBqPeExtjd4TiAWW1KedOsRLQ1gjg/
ZUIRAJCzcgOM467hlbLC6oRmeRi2kRrj31peKXEnaUe+fxWcDzM2xwmfj/62PrNFtCI8bucuNjxD
mg1hzf3PF+cREqyD84JwKsfyZiqhS9iGBEUVhP5zMXvPfx9X5q1Q14SDNBi/k35slBN8IAPY/9vV
LjgTVB7x8WxYFObcJ0VxK42ezZCm5PpBDsQDrRdsEbh1q7q9Px5hTjnqMev2wm7cHGY/CHbdKks7
MQWZ4YTrh+Gn93aMdr6sqM8nyNMf94rEyzIXpXz7BOK3ul8eTBtTZSdl5Dzzksd3mLt9YRxSyGxw
giBC8lwdnNGfs8Q/EUDdA/P3WpeJbVrxYL85V26VBt3NCr+UoCfPGYy/GiVxJtuRNr445DRGyuSa
/8bX58Wjiwkar8iD/j/WzCILg5aatSG2vx8TV2NKFdQ40jwhjkYl538QZr92f/ix8Cx4Gi5wMV62
myJUGyakA6qoeQpoeX+H5U6wl6a4+60VSimJzdK/tZ1repJ0MtdUl5eyso2e1AtWu79JiXR1az2o
xQ7h1YZZnvYS0Lh+mvhtm+Jq4JVxfeZmgQi1ZqjVi6GOHxiaShloU6OJKFHJuNc+iTSSqoxk9wCZ
lDsJBBdyAZq82OWPrSq2SkHVzwuzY+7Zz+VGNARTz4ojYSWKHPO45rh51MnJ5hIgy0y79D9f5jkY
64cFpmSNHjRnPR5z4UjRN/a8+K2FLYEu3uhBWjD2J3SndEnGThQLR5Ipx6sNGy7hBrZkENqXsGPg
u6s3kCTHqc+1uowsDZu/es7JdMpuxULnMZnMdLA2/2a5O/GEO5TOxB81XltUP125YLaTIcrxthrS
RwB1MqIuoj42BqQ1fDeyEjFWYazXGwKJNueRB9yZQZuuH1lZRQli4DLkGLD3bIFP8SdgS4znlQH6
YKGpAqSHvAo0Q1K9ikJDjXqTFB5K25vXuNmXK+PRhRUDoqU8taygbRCKAos/No2LkeDOaWLQIlZE
nvar/OZMjn4VbM32fU5GNzcSF6VM8aoDEfQLOLUpW4zoUdvh0NmIXBQuEA0ujtXsgnr6NJebXaLP
bLKAC0go/M5IjKawGOH9OsCuXkLlSHsWUYfOZa1fT+17u5CMNPrptarYNqhxLn4Shm0zMzkziWQI
6n0CfSKRrIJaVBxqUVJnSSrti35uoyx3ciTsi+PQc1pFUhBI8ofH5rxN7fgc/lQd3IFc5x/fc1Ht
bvmrQgwj2O5oL6Qx/S+YRCsuIK1S79hWsAUQ5bsEwhwgnRjbtJgrhoA1J5i0sr3+NdQ5WPj+L6Ii
kY4+Ws1mxqgu3YUSIsao/Cb67nBmGoRamNPQhIXZlsNOB44i4J1XxdVBPByYEDnXR4K4ByjYdGWn
fT1AUh4ALkMr32HwLyq7ywwQhJfSPt2BUI/tquCdm45/iUjGZ+HarISlWzVYGoty1j04e2sy99oW
sOk3DccPbz30RQOUh6pGLBsl+8AJT9+UTqpoqA9cjR1MfUtqUPqSPmuWU4b/gw6WsnWZnLjJvktj
sF5CNemhXjIjpqHxGaQI3sSphPNprFA9kSjUwyVCWBWAzVVTvjm2QutvvhTuMYSkdCTzmpmgNp0L
XM2wsKF8/t2EiJDyuvzdggg6Vxtp41oP3SqZ4athkSh/KIa7Prmhs6yUX424Ei18YPmXNcIksiql
gflj4PLi44kMlICI07XuBlbgaZfsR4hoUqg22FG1/ejJV/9dVYflbqCAoVDube3qd96ZkXgnLhue
DGrwGt7olMi25zfeQucHq+hAgbu75tnMBfTGzYPC8H5/4yp7iRH11Qmf2dFiBUWu8k/leMAgEkX6
SMEyF29+2Z2F71CQ91gEEchebdPcgDOjkl8W9YEKXpMVgWmIa33Bi98qtknlVapEeteAgIYOSICY
ewfiFAtMw0iQsLXlRV6Hb9UKBLHM9k3+4TZcyH2l/LrUDRwB99eRkVMHe3nN/1TNpbKPjpVLvktQ
yzWC0Dlq76e3ooOkBcJs/PEXgsXFlq4wwn5V2Sxbp8WR0apgmNR+a9otaNDpbX8ubXOv7+ubSNkT
d1E6Zo7k/FYzNwW0+8FPBSflntq6fsmOYkOuMAx0e/etMrbX6vjI0ow1lhZX6xHhOCCu98cGg3eI
yVQsL+5Bv/LCKz1YpUhsW9XJ3utTiicex0tyfA3QEL21oKMT/jmH+NBqp3YjALe7GsEcSM4/ufPr
/K9/Ly04pDk4KPRIdiWwgtP2ygzjuF2Hp7yUcurNegkq4xBbOGVFUBNHZqvP6rfKS7kKGrShPCX7
xFwxtZguCNyAhDOAf005QNX/ZOezm9O6IPbNlvWdNhnHq/LAxKJV9DCZ9jnE9MONM8D2L0N/wW5B
iSS2oTmKGo0N+ZU4TpsKZ8c0rOf88pgJoC8WVmIMZNWPuX3/MnHKfDed3zpE/kLH2cZ5t3K5RxrO
3vj3Z09XJcULMDKTmtvbZDwMSxL23sop9hDc8uZ3TVwQFytykfcUo+bhvMwD1O0BXOIVfMDIEmXL
BaDcCqF6dcr+jR4gdJHCVm0m7De44jok0zaVIRyn+R0nGBzHaEz+K0H2CB0TwN5xLCGi/O+2t5b6
aabVyMaSpMuWpI4+wkA6uI0GQ8+BX9Z1Dx1xLtydNw4Rz4NNcFj5bmoJ/SQ65UlCafCl1yC2RYHW
gaM/mNE14MYZlrBv21sZKCRS7zDGi5UTpSx78RhNwoPxl2OkhOiVWkh1nptE81FvjTYdTx+hCBAh
N8Mxh5BWlcRwGzKwzwgV8EJRQcwJekfHCHDdp03TXi0xdKgL6lkZzhz/tVRUnA+bp7lYSy/n6Gbm
eNFK9DOptV8Y27Z2M2FqUugPle4Q2m7kBJNUvDvgRIkaqhMMKdzZtEVP7uCoNmKn4Ytc92vrZ9CC
DGhCka+h74EBJU04UvuHGbLkbI5h71C191z0JPwbChlhrh7On/m4ntU8b5g0mGwWHw4S29TJdmM7
8DyuuobzY/5SZDRVWM2W67aW5D+uIPDGMDFVWzlzw9sEbBoMMTDZZBgP403+811qaV+f4b6vCBqr
hJd59FRXJm+EjIMApSJfnBjR0rD4sJ0WuHpOzCn9pHS8cpdFCyf4KPCr3+QYpI0oedJ8aYSt02Dh
W/Wd67l6vqhBemwoKnHVXE7trxK3L3cHlDvO5eOR4+MS0rSYTgyBxs4sRgs+JYRlT0CS+hYDkEp0
i+qUnWfHGwo8CY+ks2vHFg6vV/PSz9Dt9egeqxw9ggWxErkZggC6R84Tza5xvgmerTz8VT0GLJ21
64WnzKLCQixadsOke1F9xhEiY7V3UzdU9+6D/w3Hk3MeR1M39gRZvCyUTQkBaB4hDK3xWBCYeO2D
HKvaVkBMec7ipTd1629hhKw1wiuunXZw2YHFx2S7uB5MUy5s+PDKy3JR0iJ2PEFPFQmvEjAziWEm
vvKGhKYFdKfceB4JKpNTNLs7CdkVdlNPfZerhZEwoWRjMV0SUpJEtXpraeqxQuR2pEsdu+22MrPE
/4xRfby0P/qc2tPNVFy+YcppPblhqktw0Gu8E/EITdLsAwWC6C1zXq9HlfZMGPCfICNYvlrklfhA
wrHPaHHQ7Zs5kHIqDVgnjB8nxRf+uOO5ajLLXDgJvMCtGDXgUUjm7dMNA/XHvxlqBNUxtuy9066F
uV0cWX1wREBDg6Tn9DF7Pc3DEyyD9OmRr/G9piU9boTrcue7Q0uH25xKufBA84WhTuM/d0d2YM8m
44TakCs5eAEuW1ycW1bpezPCOQE2A9hoR3C1CbgC0eSZ0X+UXzo2GUFotMYwXcjraBkJjlXpQGRf
pphek5idRRbEHx7Dwbv5wG+VypUg4YoLi+/gZT57vF7d5rBa2kyBbUsTrGzYXDdMP30R0AL2q7wf
aPkf7MxlxnHrGZwXapiHUvlKRRZlv9IVEMA85uIvCd8n8w2XyKyAISCz1B0kfgfSq5tSwHhRo2YL
WUjLuetncsWOpirjaA8OlCdlNmdUFlcU3shOVNcE9AQ9FzWSNszJQPfvl0UZrB9bHEUgV/erNijr
VBuktqVYbhs2iAXwpbniNFvHthlVgbqOJN5ulVeMZyJYqMdck4/Xh/CA6uzIrF1tHROI2JfI7x+X
Em7Q98MUWgERz34i5EmRDtDiDd8t5gZh1lxkkIQaGU1F5R3iEMhwkis+tQzZGgzdEY1mpuMqzewK
/1byJeMLmGuX8TwHLXU3vhdQBnLXK+3FW+Qo6zMnFKSfZPYYLswmnbe6evCqsE0Y1fMDtG5f4Khl
AUvg6uaGZXQqXA9zjIxgm59jf4Ot/ketBNGlb5WsOUP/Dcl/zrNpfht+xJ4RKYbBtMhcY9kQdmWz
wGSww79LsxXjlDBuOyyYK0HCeHfZoNWZOSm6kaCFwxYEB1K7/z9o6fr/ECAFKU65eXKH+KU1ZT1k
eJNZqj98kYZl0jxKkwbXvhrlg8QyAWNTwzhQhjZ1SPXEpE6A8T8f0QsRjgImeYaszxTPF76NPUwZ
WlzV1Y7jS4IOUlwLZdkcOmIrNgGpmpySF9yXvHqXEGXkgx8UkQJ8Co4jjUbpLtpuQIu4jsfFgWEb
SRP6UOxXn0X7WOz44rjC+kylpypn2dHGSq3JHRffRDj8JHdA7sxfpXFWLidv6J5c4G1w5kk02LlI
rmGdrYbxjSuIFVVMUDfMhBj/PV4ZNEowbqzisaEzKiPjnCnQDGJpzzym2oW9nuVcU5ON/r+wT3fC
SQDaRgLvYrrZF0nad6eHEuS/HcazA4RN554Pbg41aZCRpV9E9gzXveCssXcxkRNZ4wPx+HtZwm9c
vXFvPUmj1ubVneyglUNCdNju50XgVrC2n05ZBBcjs5cBjorMhT+YQyQ5AZQPJlMTKzqHDYO7FDAK
SZ9K89h1gXq/u+LXVCfUsuHE8FhIwmopJ2pA+PZe/KJVMUzp36IMXitQyM4u1W7eRd2/niOztP+J
19HDLpz9H6540zvZygg0Lm4BO7iBQKyXA90NQGb71rT/bidVhaYqY26EXCf5CJv8fCJ9OS8KWqll
foQRanqVmcDMvQtqFpASLRAPch5lVUbWv0cb94w7Bwfp7ImFcXYqySQnVOuJcy7d+OPpsuSsFDqN
/7rrqteZ8QSpmA+Mvwec7cUy2uJZs47nrPEu25A8mMyKePUuWMc1bnZTXoCtDFzjc/ocH7aGTL2M
FMPywtrkUkqlqrZKJtZhN4w5xWgI23+qne+uuqns5nG6A5y2T+y9jT4JGai4iVZ7ecVa5RgHfsAi
ZYQVldSyZEtuCljBU/X7ANS3tkaxbpZguHMNeQouls4hDjPXsjbfNo0w0i7jLt4+f4fVNLuxkrAx
B+fkoYRX/yjMi9DHSaO7tiIUURQ7xSwQ5khFRHX+Uo4EQvxWkSxgu0gPwKgz8OiRGJIVPxlw0g+x
SKjg+FzMqXndjZ3DrLwpI9C0KhzVth8XAdZL0UBYFR8nHhb+5t1+R+q7mHsqIci1lcsl8+/D5Xr0
n5d6uUqicWNxASofqL4w27/9JOEm49cCqUDoBYv0dK/hWdte2ZXf6aDVZTIZHrWJxadfH1CYFQBp
v+IuYNlfImEc8YWJit7HkXjVjRc6wqCjYDn3rWahLEjCifuDSL6r4JJWJ0hIzLYGtG5HrgBSSipc
74/Rv3Mcv+sLr1leTG8i10NLOBfws82iA9MoCtjmYPPY9JGpg9HjQpbDdSteuY3apb1jtOpNQF00
ii3h7rGxBoT18S+5UkZ/368ww+hDtyPF7Iobw/aDC2V5gBcwVBMzHKSxNckEI5scRoilrHnFStsg
BIV2l+HJMbc3PHOWJGl5cb7HWthwfqBB3Lk10UZ+5SHdNQy4D4NHrCfEJtSrI3B6G55C5pNZFxGH
hNQAyY26dWSve+fx6GRYnYjBbb+QIyBOsDS1oKU0KVny3v2fpN4KqnFvt99TfZVBcyDXPCdqm/Kj
1bOk6Z3s/WdA6q1RZwGoX4ji4ncxAZIuOBoZ3hsJbLGtdYC+UMySCUHNYNauoSWRT3xMm7IocuK2
eubtuMQVejPNYc6KFHHCGUBfMLsuynWPKIsr+nXSr1+sEknjPGyTzo7ZxHYNe1pnYDFXqM+TL3cs
9lfqX57khBBLGKveQAV7DuQCgU+ZTlsbMpE3FwqZFy2uQZJsgEi6kWB1l21h1lpQqvl+4pe9zIXQ
Qu8ZhYXolD7vRhDl9uIGRZJstOD4LrFj+oLj370FaFl7dPlD0a9qF4Wasui1XA95XMylX1QyRhNI
NDNqR5a+qRu5LZXL8lJC4BjVUv63pyj72t9L10kkIC6ELnhZxu8ZI48XxZjGg3SNjV0ErYsvpr36
HsAx8kAEhRcKwzFC9Xhwxt7XRc98z13xEYaXnL2V/S4oH1tUfQcdBJxesphwruUHQAOhP5qujoc1
b+aWbzvtTE8a0mzYOUuzOZOty0JLnFan6ZkQKmDhRAklPwYuvTkpgOo87qlcJRAHh+/r0oEpLe5j
5ra3IRWWqtK7LURq0c8MMcddyrb2wZFFElgvG+BxtDZSnk2aP4fve3PJIXTLsQRaiOISCejKF1jr
OJYoWhV4vSdtJyHyCbxhlkC/Th9FF1UyXZmynMcE3J0Q02+m3pRm7hyswlH6zWMhkr/ifdqLHlsx
5yXoiGcWhnF+JaBFlMrf7JJ2qoEC1c/JFwm3Omjow/V3Z101/e9l73c+z80dh3gFAtGfHKDh9dtW
0DnI7ukeudrS4zfRy4AdWeK6A1p74c+q7xaoSqB+cRAZH/vLx2V3NYRN3CKNhd4SvHYCECiVrCW1
DbBgWfj3bhQJFkrfD8DsWd+GM3FzIIbCh043hjuK5+cHJYs5CVOPGb76kPFms1CQ9vwU8ZOCrnFy
JHGZT4zjPyhNKraJe9EdeJ1ZEoBXYyZtlFceLJO3cOvq4mu4V7xEFEQ5yqPKT3C+E3aRbZzicGpk
efnacmDFZcUgBYT7E+yRTyzB2ctJS76rc8Z//oX16GixEGqPt5d236yjef6QSj7zrwteynukwyOI
lwBRfTYEkn7p8BMaCq4fUU6YyoVZrkb24poQdPFQHEHghH81AI0dX5xY/Hme3LLV6xHVTAuwQHWp
SUWNGlijNWrJMnwhvngQ/wSewkKe417xQho11z5YpxhBBBo0ToA8Y1dJuFknze3kRVryB130YZ6k
qGvhq1CNJK0Ki8dBlRJ3zkLu8wlA6AMm4kF3T2jTTP20GSXQ6UELO1DETWV1jjxMG6yUGUJpingi
fs5rUFkC5K51NTv+5Iumgd9EoROnXUJGTelgpYxUVkW/4v2FbW0e35TALWibI3l1ZsspUxD0yRWS
1DjzuCSvfzvdREBbHlMoTZZzwtJmWagob1WRxd9ju6zUaS7XyUvtA6E/jZkFJuhLvcrjvzvatiWj
tqYnjTyuQHYs4jWx78KXS5VYb2yJ8ZSZ2OxixhINyZG0N6ZsxceMI0o50ga76UZBMSjTwJ4tABYV
CXzcMj89u8MuhxzoWtlLDWz8vnn/rp1QbgfvheGyV0rXKtU5dW9AVdkDnF9zPdyq0mV6mGT8i91t
N3T0bmHaydOepV63/nl5Ubvtq+XE1jjIWxp1BVVB7ut//mddmQHPh307gBe3S1TcI5gLrg9X2KKc
ubYEROsFXbfQmuy+Uu0pIGlW4xQ8wsxnZ0M4q/BoenGbp+IGqalOjYHpWB/xDeMM8ZRc6ANjxRpB
+qsmC3VpN9UGTc3wKndRChpAaDsmrP1VlXUkv91z1VzukiVAPg6qz1vgrzAYzobmQXkvwjUcYSmL
PrhZedM0CVXvforORk8194CPLBtotUdZEEoe7Wl3KcA7FWdp1fZ2yXkClsuD6Qo1rGP6DcClAXtH
fVAcuKYEKSeJdm2m+Us7cu2vFxaErcHFKsqFbN7DIV4duLpNvUIiODKBD8rHnx3w0VAZ8grgG6wB
68ZXXYvvsBQIUdqh78lzOVKqA7yHy3A/31e9vRgsIFMEsZ1N+yakpv8Z3NpQL5Pouye1oaZlvfO3
E1/aVzvPi878HtE3JjnOtIEmaMRcqHBucFbOjSwzgHhfHTrQFwoKvD0dc09DJPNT7rQQRCeJdR+w
8shVVB9m+KSt9FvxDvXg0bL6fOIkrSg+dYBMj0G5Rjub5uKLJxPNvyO/Q/aSFWqVh4zjxSLWdK6P
HHZM8gQglZN9MFVPS3DlWQTLRt16ZCgkM+vQ2gtNarbcThaUri/u99iRWHPg+Rt2ooCyEtUVquvM
x4qMX2pxMDoRuq7HuBKQ6te/oxBuowsBvB7IKsVEYWm088vxXVKkQmN/Yop+Yvo3CrZRWC1q+2RV
TJwJDen47Mje1hpH71/kY9/0IjvdfmVVWVvKueLpRBC24Vt0hGXLUdkR7H+aLdEP3XUhFGUwtSx6
YmkEgeM6WglBn0zvXelZejPyM2FhbojHd+El4be+gnur2xuqek3qwfaQnxmGacOO5ZJN/tDX+mml
3cnYLBHXi95ijUPEElNkVnvYgA+MaO88Oi88MtbBSItakC/ol9uFVdiu2nJcovMI+Ezggb5V110C
DBtNpKD4UYNtO91CwiNb+sNibcBz2apB7vZSA/6+d1vEmfZ8P5xGhbCRvgwcezLGr5B8F3GeQmmN
0ZaJ3p4cJZbrlcnUyHpKDdokDktlUPPPaHdEQWQDJH/javXARiHhXpPKZUMWobbWQZac7IYdpwRN
qeS2MtqQJSloAIModc+amRN34QSSDpFnUVOJb6+bX+FbX7bIPMndwPeb19irY98Hzq8ci6prLPVL
03QZxraIxVoS51cxBznhvM8Na2TseML2oH+XdvM7WmdYD58b6Eznc/c7wYAoYNsfG1jIhDU7fzDk
Njk8wFEl6wM2cTcN+Cqb+FHm37G8waNoR3RwSr//SgQZ8Tz/+dcmxVhO+JivPdDeIONU5+aR9Mc0
dbC5yrEa7lsFHvUg3mFfi8o0YcJY++1ilrCDuyR9cgZtOOpG8aDDTJtnRe/KPocmv4z4D/IR3o8j
+zPYOLnQvR/cmcT13YZUMuAOIy962Pn6DXjXXs1oFKoSiekHOCMnCMXqHDzfOSmHdSuaUtqQmO8R
h3xH0LKrBPY42MeSr8ePZ5rbIx5UqZbvXvLQ3DWk+W940vleIjiDvNq9JD2qjKt4sCJwqmmI7qk0
iAb+MjCe+XCuR3Def1s1bDP9cymuSdVjiExLfMOe06glhmmm3jS8soHRzfR6gQEPCsbRc3qMnGuT
v/7ZvnfbkMWLsaHpqoE9MtSf+bDrUUoqRX7e3wj/nadGf8pdz5v5D9moJaIackUffZDsFCs+55mE
Yk1vB2DIyfy0deQsIKFkDES3umqFpGkg0sqlCUfbfu8g8X9CmIVmoHiVD3ZHKCo9ZXBvmvo36Q7u
NGZxvwj0ERc1+hztI+lwO+qbDHLF7mdjn7AmGI8JWoTnC/ot4QnSBb/89hAnq+K+ZCfU3kaWi0XS
rqzT6IPToIsZRrz80JCk7CdvaZq003jKF9op1CxfJqEIxzHD4GAPlyHwljUeg8h+nEodU5HDm/kH
c8k7TBxn0dHitE9LTa5AerFudEpY4lLHpxahjBRQ8Wmyef2FZ+waRdJv16FHF0ZkyRgx0p+Pg2H8
kxairG0J+lR22nt1XKTAz+c8kc3FZVMH7oabdsP0iKin+pojSm8hvMkOXcsq1tYYssaacVEGhEyl
iFxiTs7afoKpNUEfUcKQT0BrVojcHQdTMWeQbQNSAUEpivo06zbe20jLWr87F1kRwkROALZJa91W
/kyd59LHjKuYQk1aVy/fklLO6adIpAcVnUFOEyyefB/uFcFlJa/d6tFi5sKYTFlJjPlI3+q8e68b
2V2QobZjLHcGNMwqTwoN5XJe90HbcAQh2tGC/WvTZ05jQyMDmXKIx5iawK4755hGo3jYvaY2VJ31
iLyvYR4V6y5oINqhwI5U/wBsxlKOy/7V+VS7Pmr7jRONlgMBS1RUFIinumOORvduDTU+Rj0rlWsK
cj+s08V++V1qb5yj0ApCAoq6Gv2Yi7WrnASkQwH4pCcx/C0r68msPIyEwcvoXU7E3DtNlFT3dVV+
qPmvj/v66IhQBEczMrxz5K6+UgE14TRuJckkEfPZMkkARETNl3pKsqfe78OGcIGQ6DWWN+HBzbqg
qvKE03GLTrJCVIKCei9eqW4rQjRZBgkBY5MOosaMCMeYQ6MBW6XCe8zNCfQDoBrdIItjhrjRKOSR
cTawFz0jk3C26J0PdFshUoYtrlhrEBTquJncaxTVJbxhbCanoDP4D5dm2cfOVD6sYxTOCf0Cv6RO
gBwXTfeaXY0L8vk/1bzqIVr9NFVn+sXCwD2dp1PGvH02ybOAUGSycGECySvgdHNSOlVPZRY8GMHE
CuAjKJA90Lsu+kvPY2hzQxldrniPEOcAL6R/wb5BOYUio5gIspenzOhsjfULxd9jF7Z/2TbzgmM4
I5AoP6Yrh14ZJ9mta7YAutVwLyVsW8cuQQk0RVbrvjhEsYUMj7Ses80u0DGXuKSJcecQib6fbUHr
rpat1ptmqtpbnQqP9ERge4I/KqcFM9Rm7etMf7H4rVqni5UZyv8wNVlzFYbB/lru5k0/sKqJ6OwS
sgcW2lXFEqjX6cZ5iyAhv3aP1PGbd1Y7EIofxTmLj85+SgtbcPdqPzmacvU6qcb4RPz3nIvBgamO
j6XYQ0s5pkGn9vGW/bSDf6Z+eZ/EqHiagSgPbWw9RXQchc7siVNNHi0D+NNNatw3fdimZaeQX1jU
CQSQqvOHucDAN04o3YN5UhK1Nl1m06f2kSCIT1eu8Dit2UX7WowCI6ycZJaypBwUfe1ULgliij2h
LW55S2p3F9Gp7Mn1ofPjLUOIRqGsEOqNxhjQW8k+XMkJOkBpNny27NeY+vkSYIFr+d8AqaxGCXTd
exqLFL4LE/wKBUfRiPVM+nHlCt/m2lPPSqedEWSSUU+9BCtLaYLhB4mzT82NJbl5UBFu8VQO2BGW
0KhHgxbPbGh7u14cgqe9rQPR2LjEE0aUBPGRxrHj6vynhxll20QVsm3EhwFLxpEf0Fb0CVTqkcLG
gxJctAICcrFTgaNqLSB2EpE6hRO/8WvvPUzILBZRGDTQU9L7vTfAqPjBby0/8+WphbsLxn8v2L4a
Zly1L0X6G6ho/hh01u24nlBdM48DglxW/dEj7jKUJ9b/3Q8U0mc1B9OXXRK9xKpCzkak5w+N/Qp3
dk5QRUfmdADUnCKF/bdem0p+UutSCNV1K2ujOGTCO3ABboz7ZgjPKaSSalTWcbGgT33IjoMy4LDV
H5NbEqz7M2JwV9UD7JdDx9feL6ek6fsk2j6Y/1jg7sjp+BVcgJ/ZB9/5gCdgM3u51jDgtCwnvmYb
MLowJ1W9GNa+XmsGgsYMprkW5tKPNeFWA1GibHDcPNWIcE1d+niwOrRFvzfkrE0SqxpHCJv14PXR
7u7B0sqNw96Q2FdSdmJRXIweyTNaXX/p7O0IgqArckxbVqbFqubL86wOAdQ4pWbmu3As1ofIBLOG
OxA5lpGC01QihYo5FXw82vgLYs046WOZyXY2Vi4J0FjgTN0UMfw72AllYExPsM7K9LrFCBT0IPO2
JjlycIA77juxQzj4pxPviIvCyNZ0q0NbB5spdMU+/3BVRGgoREPiU8+/dVosDM7tpq+Z7p7J15Ev
7T0x97wWrVmxHa7OWShzo0SSTUVOCW5qhQVzon6faZCipGRK2eZRAV0rdQuWAmy3Cc6YihX3frSx
YxrxDimlVs175IidMJd2HjiIPFss5mZ0FjvP/uPSlgUsQuwyqE9xMO1B5TZbzGKhICWbO8DFrgKw
2iJaC3toRja3dmsef6VgdxlpJL8d23UQqr81xISVrPJGBVbxUUkDTvFOhTMzRKs/rzBQ1UDtuD//
MTfHuqj2ap62C1HSx5WlW9njDIfyUMvh5ZihcBhsEAM1zH9BfnmgO/FSGx1e5dUbLqiudlD2qDaN
VumM8bp12beTmWf6j8AUsC/6cv7EXqlgCezFPAEbVQ1nYueCXAAdxcGwi6qqePLDtITj8jsFSBWZ
DLuuEYuQ86LauDCA8mprC0xDdq1+//TMmXTDTfC1b6+Q3UcD32LeAaCC6RQtsUIvk1n7AS/w+TLp
gq0DtyJdIMlPYCs8kcwDozQdnvZxMS6zkNalIssFYxWCz6ANnGyWR37yebDaUx/D8EuMyKufkxyz
SDjmb1FuUPD6p6eqdAYfkHVU3U+J1HNirWxPB4uRMAtI2Bzj91ChfwKrK/0G7j6gbGR6olkLzKAs
uvLLuug6coVLyjo3mbLydFe6Qeu3K03pzm1qFGcPTPE2JRrfkH3Gf9s/dvajsRUIINdgfKZnMaNH
gT7Ss2bgFt12k3Mo40x8MMfVmnoTTMOVB5bQt/1aaJ0NrCAnefiUAVPlwD0eQcqHGDBZEciUhRxG
Lkr3nrmCXibDBrQufcGLJNDkbYWCwjUbC1CirzJRWZIPjl75e8T4NdudFCRTKv919fCiNQTrn+Xg
LoMQuM3N0OONcATSI+S14wGW+HJu1lkelT/+rAXRh/TrvnG/impAGQGKb7iaEpur7g6PgqL0bkY+
Ugi4fDvF5JB5fKNSS53A8ZL4R7jE3Pu/qOgwt3R7LwvdPNjYqn8aKGKhgM7Lluon/ppUQxThNGF/
EbpS+KhtaCKAz2csrAeeOGZ4hdsAwYYSUKqjgvdr2z/jNtAVRBPJkr3H7V5tPVS8YgKJb2Qb6E+/
zJRtmm4IZp1C8BNxmdLRUwC/5baLcdLewTOWEw/On7C9eg/p5e7jBtvsDwoOGTh2li/venJTKw3M
UA1PE/gFThnVUcqrgl5dtbR0zScrKJZ0OMt3k9Hmcvk5ZZAqh06QjRdXmW/sO5Zb7eL5G6mJPKiq
pr50kELZY4q7g2ffcGO23SSsNMVNvcbLTD3HPB0KUuWr+ks+oUGy7PqnOJ4PWUok/MS2LRDKlwPG
7eFWCUN6TUdmAS0Ipj9JHv56yiNUfuAJE2ZWfWtDwUMTY/OH7yGbhFUTySuXa7KaC56OuQSy8wP1
1qKVAj+ZeGqbgNMamyJbEyri20hJZN5uI/WAEf7PZUzrd+Ll/ICbkJTLOOtpHZNCeiacvcHGIi/T
7+JQSSK3tJ7OdP60SLUXjMJICgmO3/Bj/23sh+efLkMVhExiHOEbu/cIq+WjBIChQC6+IFAIByRr
Yp9d1/Dct0kMtBiZ4XaQCO8CdtTWCsXxQG78a5eRiG5VkxxuXFQJupzZJCdx/WxLjjn6+l0AZFBa
sq/Ilb2KkwqXO3+9/GBcVdWfDSsyUftl6pMjc7qzL6tdmtrQlLjRqs4m+B5yDzLTRu35W/JhzfMS
zLnLzjwWu4222rHxlV/ScJW9XMFoRflSzuYRsLa7KQh7+R+qwGkVSml272Mg4UvUNLl7NpfNQgOI
CBKlGZuUIp2a0oV6G01r+Y+oOwsgQzOPlZ+PrzIeN8hBARbor8o9pUSDNLKHOxGCcp0fEJ/4LvJq
8FSc2psIrs28Jmd+OHWyyHY1cCt8b8tEyerhnXq5+DqWEiT81uYKhBp/wSnsxAda6xqB1jZWicME
UKRUjZU/YX8v5w5QjAHFCS3pUIyTNEh8P6t8I2UZXPyAcX3IY37M1ZrbfHSje4X8X/+gnM5NRKjc
X72bbaHs7Z6UdTUc052WefKyqBTyU+i8OZGzMzSIzH1VORuX0Tm0yaiHLWllM9EuHnCH1U4A3u7c
DcZ+SjFit+E2kG0YwZrOTyUKyjRQrEO2EVKGKFu/f5Rrc+iYNgs7tMPRj5RD9LoyX76spyqbCmG7
Xj3Zes6QOZ5hkqLwWmT7hz/W8jQs7zN8JpVl5LQUL8B2JyHSiKzq1zLATQRZWcS3B8/0OEvFjFKm
2omqatWENzzh8l6m+w+rPCt6T9nHddfAhqWht3bW7QkuRBT7DHLpj2dDUDVA4W2R4oYlNV5eMFks
12XO/mjNGeZ1eLvoBlTQmLVm+v+49Mk2whMfVGyKGQH2w78abc2hE4IGQH+Y7jEOxe8BgbFXegS7
q6qEpqREjdN/uFOySfT384tgD/VzjQAuC40fey+NzRPcKa1RdnLqvBzhfbTHNDMLXpmETd8Zl8ld
djkgEjMngmM0uMdQNd1p3GyNKKkUPu6UKQrv4tn2w3+LO5uShtf1PIu6m2mczOkr7PU7ZD8LhKEE
xoLJ34ILeRYtybIQioWwdEYToPCaYJEQZ3J5x+HfB17xc1JAdAzgxQgSIlBO9JAYLj7vFfJr5q24
1TXzY/kjHmjwfuzxBI+PUTmVyquJcDCLvnT4EGBX7frzGUEm9lRU37RxZyZspVvPBtzBAbUq6dIb
vSE+r8G/hW9AviH506YYXo2epxEkqI4fWO9Nuah+aRPNZVLYRckIffAUsqIbmRSQWGGcHZtyveJe
DhqqVL8eMCJfyqvrHT8PRtFgc5TqEHdDZUueLZPKNxy8NNLDKtAKtkXhYvwJh7i0w5AGzOxrc7RC
ByypFRXW/vHTZWtPO1FDLmYcNy/MMRwqsT0U0gtycDGh3lWW8bE+7nQzTGD4XIJ5b0pcbTN26Rzg
jAYOHHfK6D7IePPC7gESgPcXgfiHpnGRc/+M+xoF26TMyN9xMAYH8gDdV19nW7+PXhAV61hlpixm
ePyZGoIFspT6RPpbkwdQStmfsHyfsX38mxVVw49fnpje/cHfGb945p/NunI+J5Cd4mllJeLcRqG8
HEkB87E0EZDYGtpnncENdjjvN2A4RzAVYmjg0SMQ0d3qrlb2npjdE8o4VVbTZ39qz9LQPieIGCCu
lfIv6fBNWOAwq2J6G6XnPx0flJDWAlKMje4sLE4p50XjNZEW04yAOiZNMSpsP2DR0FRRB/0GLxI2
c23gkCO45U0HmIiD7vgUVvm15X74pepwivyAcnh1xdCfadER6D88JJt9seLKUQo36zlE6IlvJ83o
XYkz/rjv+3eQ+tSic1TUuJctTpB6P4tOS9AgrVo8fFXwXZKK9Jsdac0POfZ9fGs8PqXFFXxlqxlQ
Gk6pUBtOHIwX1EQ4MVK5omTYmAAwdhwiJni0hjjaaaKHABHFl8AG/fxY6ioOvyAXFU9ALBI1N3wY
acCOuzeeCmRO9arFpIGi/w6HelWygyoIvqJQDipvjxmomkwEMzzOWI13Mhw9jJ7A9GAK6HkNuMpN
DSsmbgEIgW7qwT4X9CGHiCRsbO3+XXPwmtXQ8vJdJKfmu1yyFW06J34iGpyFE2+GfzmmpoDt4KhB
aOlRM/+qW5H+HaQQ9ExAnWn5nz9FXdRL1MPQxQSIke0mlZgereXLQXJn1PuMhH5U6sa4zyuTOsJe
b/jfJiCrMEGPolWIh0nAnDRegMgsnu/CJjk7+4xW+INMiWCnTv1VzybB3UnTXKV85R5JDPmM+TCU
gon7EeY5UodUVmbvrTYo0iIQtTLN1HaGisnBlp/9sntJ1wYqTh6GlFgetD94Dtwp3J91XihCyAQc
HjpYiPc3fZAWdslbzo/fTXXajOdM2FUi2xu26zUMWix925UrUlkv7U5gwGPojKRkvSJlW5xnxbgq
/8BZ66+rO1DVDN2ZUiqQK5JxqQ1NGU8KsH6AjJl+TCPASPPXoRzyUytDxAu7DXnwjoogRZIGUHRH
vJuzaHY106t/jWvFkqdP3pZKthZbHFSDEYQfI6N5CGgyX/SKfiavZ6HmuSsqS1esOBCihfDh7yTs
ki8cKgfNjPlZZ3/uwYNkw6gvEknTbgSmbxGKDEqs2t6AcpN+GoWFufpLX4EqouZzJRc479sQs9oN
e4q6WkLwDKbpdFeDfjBowQkGcyGdS9SXpMSNs4BqNbh5/atie+d1q1NKZyOPYEVk/5S1gCqZSCwJ
w30Kz0gaJmzU8Pssuhq65qo5VdWCZaF5FbT2Yw5XmpQbclMXDKJwFn+JoGb4kfta0jTPpCqMC9NS
0uvNrFMeLHpiH2RLR+F2AKJu1zTiUAazayb6AhazyqhOEnm1tL98Aqu77acDg6MLaP9J0ZgbyFBu
K/QgxAN3/fOovOhf7O2lY6638YtATAhe7kv+zmeyqyksgd62KDhDASQrfSnKFsUTkX7cb/fQRIbV
AMfK25t0rqiQZkk9X6h2VzE/6vVN2yhYTYxZehgLryjRzzAiXJN+lRKMYQUAvb0rOxk60OqMx0gh
H3OB7E+dPxhTzG8mt6Y4VgrDSZBiQkQWZ6mwkaZM2h+FDU/ol9zKzMUO0cSHNOavkUr8RRv2xvHs
oSIn5kimZyVLm58+5MHojiv4z0gnbgVsPddMrfuvA04MiwvUFFfRdEQ5KE5kyn/ixFlHF8xuiAUe
pbAw+NxkHvBU+8kV8S+2nszJqe+NuyaNvsPuQb1T6DKv0+1zxjTXR4VuBbrBO687ULruZ5ELqA0r
5+yx2/UdavlB6o3gmw5YJszKQTldPMQlSIIZPKny318fBg7+LFoq8QKqXsrcRqCobZ/XLp0g6hut
z9du6afVnkANUSMC/BKbre5Znv3Fw2+09bCQiqHTjg2mrcXmqc5GMpcE8+BJjoNTk9ldY3xvwniQ
+auCH4XnMvfPcjO/yvAOdM5+CsxAZo8nLiRWFQIPwlMHoTj5Qrc9vasOTlrQzx1LO2JgeIZJAzDj
6+VmALJNEu8jy86q3JKyjSAfyu8IYj7pORaCid6ruTTbKwHgOLnM1uwHOwKo6pirLc34X17sgney
myQMnL4YPM4q0j5hBwXrg+YsTZRtG3xlJqfYfzFAYzeZ6vOtK0BoU+z6JnrS67ZCzU5u3IA49EvY
SP6sCEwbfWzs5sDCvqEwilhEVOMqw/WExiJddLo0Vw5ZCs0JobfIiUrIcRxGrMpDxyTLyZiyHOiu
w+aRYSCKXZyE5kChJs7ZRdLWvRe7o8VbzGOZ9O3tWE3jEzMcheexY+rgEAcdbtjMqEmo4dN6ZLBp
Rljkq1kf5efgYF2K292EbeSPkVijbSB9pJnAvTKdlTqmVraBxZGPlOLlXDeVimu8lAqEQKYU1cJg
z0o4qoNuiM53Aa2x/lqangKU8WLyejGC3H10KlurXR91VVO0pZg8ovNtp1Jz8BCogphHyjXv2OZB
9vj4LHVzSdUQanQz6AwZEl5KoTEI8udUYE+v8c98zL4RTVRVZFfyYN6Erm9OJsi9bI2eS00f8ny7
J9p+PK9bRHhFrZu/R2dskJHjqTETkNLCaUlg4CihtjbECNqqOd84bSKIl8AZH4jSVZRSFXERue6k
HeazGJW0+eqwGUlnS6N4gG7uC+skhjnLYEqn14Gb8Rgch2Qb1es9G0EYSHSQg4hsPfjuSsNw+sOf
zY8ki3SFELsMGn7Leei/wvPf2ctnk1WKuTEOTJP5YA9Cr0eqNqARMq+OGOb2HaIIsI15gDEWNCST
A712NVNoDQjeQc3Qb99NaEoB44nA04EPZjAt1/UhuofXBs1ifp9fanzz9CzeZ8uPTRFUUAwR8aFq
kI1F+LYyEwL7vnh13n0G29Erix6SC8W0H05XCnlOzgB/QwtqiL5HJx8Fn0uUy7/R75WGs9OkWsZS
nd5VPAv82nqw6fyQphIphoS6txqPsPvVHaGTXWMPRhGf5dDScqRiuGC3Yx2J3U2pmo/i03A3la+U
mMgEOnakpR9k13RRt5OdWt0etzYSoFuWpcT6XKXL+4ridM13U5ZU6o5rBQxyoVlPCbYFABWHQfcL
vosX9A20wEPZYlf/eOviMA9po8k5vgC+f6Fiz8/fvULIX4D15xEmrBpFtyrep7tcn8HlrIzwSAJ0
ILL8b8gQFXWcq/pyX5eYO++Ly1ZjGfLL2FxkSNDegQlH7gfK/xNugS57OXF8/muCdmGDM0rkQ/7Y
l2JDLt6vUF45fGODLTv3BoCkiItm2iMCvnAe78bOcUSqOP4BzkqdZLG4xik8XBIWizQu/SwNDfk1
Nne6sKHzdO0WJfQx0MzCOMsnXaTtg3yIB1VgvRghxdR7XE+SVjkTYYiM+N9hxWmrgNVCcA0jVNWA
175uwYfUgJ/XedEDKbeH85CZ8mOL4Z/p0N6rTc2xNe5/RZZvT7OBDEepJZyojBiCzbB7bmH5nFnX
wH8Q4Q5Hj7pKujNAfv8Ljc9113ZlpYmufYcCUFjQ26z5m23nTY2HDdy331LYA3Qk1K1VrYMMOgiv
JLVkunK5c0zsq24PX/+VujIaZvrtElWxCpdPFadQ8n+7c/gatceT5L0I6YZvG9MZOAqJLQEzuWes
6pwJd6q5QzRBjAxTuzjmCInmNPOcW+1P8g/5G82TXyE22hxowFIth4J9QfkyRs1nYdsMVTCFThp/
uBxbYxJPHJZNDNehNh5EBPMowbewTHToVOOMUMB8HVsMTp0VX0FHs34n8OXwrqRhvAzJ9fw0Ady5
l4Ba0vENgQ4LEM8tqGCSYFETyMyAum2myCy6xDmVkfX1ik7Uv6ywaqu5p6GYgEoIGN4jekZv4q/1
ecFwdQLBusDqzsikYeq8Er5dJmq7mkovHdY1YA+ZvSUOB4dm8OScp1K44rJSOVnKRHa623WTAnvL
7ZSekwsrrIRY9uhOfuQuWqzXjO3xUamhZKXiovNBm/0y4NIe+nQYedVBcR2AASvGbYiUCZbEupur
ZGTEQCJBaO7vEr1qf0U8+HAmVtsrvmfNgodx9cW1Mn3LXkhvv0A+N9gdabgP3lv5l6RLvM6KuZTe
+bcKkKWvrWc2L1wPXLXx+RfwtoNfUyeI6uBssxrElxTP7yo7iLGdTNv4tNgol/LyQDLFjHsk5c1G
CXk4dIAmQ/x2BNFPwFkgf16DvvWSh0uchnSJ6/KY80pvg8xzskGdssEhkSjNvkXNTlBdmOaNT/n9
VmiOBQVFQUTT+RjeTHR8hq0wmv75y4ZvH0a6soVKLeYM2C/yy+qZqDdHriTYGon0WFaR+Dy+RizJ
5TI2Z/AaC9ux2fB1aE81NBqXbm19xiwqWELH8Uk+JIvIF9YrjZs95/Q2/oLCxhD3MwAI9G67Uk+z
h+Wq+ixfkReRxnUXqPfvbYZDo1hjmd6dhpAkvKc3b8EJQeUEoF8mdqDT9jSUgzoTZhaVx9HJH+as
eWQxp3PWvkdmvRUY56W2m4uHMleculBe1043WhJEUGyKhCYQxzVnsFDmHuACtccrn8f5ttmCHob7
tecUxigwryixy77WBVxGlll3pGoIQYicPmLQBwdVLYtmfZPj6bXh7UE3X677qzzzFQe/yPFTKGmL
bjr2AxVMJOkG0u8yIlzNHJg0YmdZdMAAig8BpxJg7/XsfBO6GDglJEuqDtsZJL2AA4MpN3pl7yHd
KQ4Uk9kt6NE9lFTi8QB7xJvCvKKLpavnN+lJkRKcnTdEm4IrpvZQQM56p/nmgLYdfD8+vhqUwGWb
xfKvYTH/v7puv9HV+IjRF0lf20tA3QE4eWnoB94R4Zg8owAvleMp9Xakc5iQ50Uv4IBPu0ZzOPe9
0+1yh0U1MX5bnovB1X2ivZVcUdB3i8rprkoeVseO/rmbVlenQiB/MyMBEp8PGIhFbEy8C+Oqlekb
w2c9PxnjgahLGFU9lDmI/YCTz8zrT41LDjuLkCxMWcYj6xWkW+Qvf8Pex1ukYdomjR55sR2qk9TO
Iw7AflRRCj7UYdWK62ylYQAnxG/KDzFoi+CeRNmkskhLylSmbSnpcoFaVmYMS1+cjbgdW6k9M9qM
XboDOk7+AlMfLquFPuQwIl8qFLoQ0IuwieJJ554DQTqT3jaDpbiq0L7SUD5uuXZAzgN4wpxdzlRz
RoAb3JeoF9y9FTENanUK09xKcO/ic+45VbFg5vBEX8G7PVLAcvVrEI7ZgXXDeYkpqSscnuu5Yq7g
uCUVnrzONeqt1QCqGMwIDO1B7HNkyXfcQkHBnDLoyup+kKg0MPKH3sAz9Mc1f6L5B2jK1U7pyHaA
Sk59l/p/pTz9wTNfqRpVqvQoEfOqk1hP3CyRV+3KBMXmcpIT0nqxaHQS+pV2D0OQMN2G248OFyby
1jRT1I7/tVX4TTOfqTTkBRX3YMOEt3gO2USVY7hEiNhNn/p8C96vKhbwSYzmuE4Zwnzon9+gPpp6
EoNzfVDYjeyE7Hq6BVSm8cZI6hJWD6jJPaArlWt7xq0SOgtDu7vUcTC06v6/6L4OlNppkxyULR03
uoz3xY7+c49L9LKvzJY+4N9DxNQZyV4Qlrzcql6ccigfUPmVl0NF9n6/Ui5JxrOQkocaESWVbvBw
3n5lDYXgaLDMbA17sw9hpk868w+q0hEC+fCUDbcs/XPMqeNvoZg1dytQLplsQgGOhEgRZ5tdoOv6
HROcxTt048dsPTZBwrsNcj95u73k7bHUKb/BDDsrjWBEQe2up+QFv+pECf7UB8tkppu7ScLEDti0
EMS8Ev4m3+2Pz8npB6dKFnbi1rqBout6dr6HqN9d1wWQ9NDMJqqu47YdgiymtWIXsoUWPpKx+5Ur
0HedR2bUVUCGJ99P7w+cgnoJqDUuiOf5fR+GsK5lnF6ZJciQ9PQrnWHmYIR9xlr3cuYEeMe0f1C7
2Syv3PCKDB1I2jfNFdtcJDYVm3qbSI86Ol9SHDGfwKTBeVNAL4B1ETNnR/y23o6q9huroyX3yAxy
0LkMGjpL+qqetlGszwcUC42ilJa3j8nMEz2qn1Eg0KdOmJI+wd4GzpM0saVCgJF5OLve8if8t+WL
FOE0niJFIDvw+M/BT6XL1lhngesAhXCFfxRGtoPENd+JO3EOaNHmn+q3TFxSrwAXAP7r761L7spH
h0TdFPjvjUiruHVNNJRN1AMUBDV/9D3o+4ne4F+go8xVwZsIVGEjJLm7xE1StBXE4n5HWW0QTpcF
8a2XC5g9Kmnm3J5RkPjjbERapmXpamZKG1DoK2pNOkaKCQx8p9ji3YK199mltzPXWm7byWJk14/T
zHPC8slC4X9p3g+DM6rVRMbJGk4mKFv/iaXAEoC7ML6B7mACf9jht1OG66RyEEZ4Cr3Q1t+sT5Te
U1d4jIHy9B9FCAdouz3mH8yPZiEARuLSgjVcrVi2Xywvyjoxv9MHBTqqlXh7S5Xrpk2/vVlACei0
GA/buFCqm5LZKJmQ8q+8zHuL15XGbNGy79wwj/HSDbkv4yy+tbt/zBZNYmhn8uT32DHjKx8hteBQ
Zy6M1shxafSs0hARxWaWy5hKf2xR38BIRjUNWJI/i/fDL5ZIfZpyD/Y+21ISomfxTEBOVr2mQy4d
IOvxmh3Na0Mk6JXtEx75aDQ3AuwbWmb8VsQUWWttCQX81nG9/5A+ZnwvQX8uN8N/L+GJRVdqnFFr
b/ZVS4rm8GenhfhxvZymDlWyd+/XTJk4sVVjZo5y8XCXltaWpSwISjmXUrZ52mYNr0a25W/kBK0f
dm8X4Ir9wpCDZM64dl79t6g+pSB3dXRSWFMW2upQe8oADepxhYFbfLHV+dbmGMc9wZkfpETcNFhz
POjXMhM+xdTpAKUgFd9+uZ7+2Zr5No5DlJrSzZkN9H57cwJOOVPH32jU05KhxftUb9Sv32p6itTl
kZVKPhA5W6VBd7UqO4sw0PZHEbeoZyKMOrjgEMqDX5+EG+f1TvbC4XJ9gkBoGHJqXUpaDt/E8CPy
KY8T9MkNcEJaE6NaO+7uGIlV5lf6YcL8D99x1diL36DUaC8vr4/ZRvY3y57BbBjMof34rpy7ESlk
7uBbrlSljIX7r3K78NnOYRC5yn0X9amWPaE8RnH/eKlOpOxOdJ6C0XJeRw5xKbKgurQnZgnxKt1V
PhiD25KAB8hT0RYv7O29kRx01zDGtmfHTBhsD3lLfnPvQFQwb/QK9x7Cu17ct6u51Sxju5lRwe8M
8SxHvv6GqJRfajpSYE/KNOUYYSoMKQXqYcCA/soEVTMRvBYBCDEERN9PJ3JBarIYRopX/B9Jp+TC
7atRRL6LqLnFwTDB+fbXGPj4cZPrVizsqW4cHHlV2/9NkfGrh34C7JWjXOS/eohJRVKBWanxAD+k
zCk+cUZCF8YWuSwhqGCnN3B02UQL/BQQw1ayyfi1Pke9O9BTj6SofVzB3rpfd2gupIAed3gNKVTu
sSOycIzg9NnAaGTUIhzgIjsVyxxyytF8MHmCHRiQLlzqeGhr4jxZOYroFGp1imizf6/8h3Evd0tw
37bTNBCfixmdZbTBIRHr5XkviSf0v5mZ0mJvolueeY1lCQxt5x8mAeRHMzrpukxRKhrjueduNMKs
k8Uocig5+2lmIC/KPagqhgZ4YRQFsSCBLYgCQ4dQJtcuqtxbIDHixJjWaaGr1ukpE28TS7GsPW1W
DuE4y89vgarbvWGk+Xb8LRVakMyaiI/bj4920ajWEaUgMz1ueoXAECGjV1I7h5O7O4O23fCexGsT
ZKOCH8QeH769B0J9LM7MFPjSnSL+WqA1YuB4kGQ6k2QRiqQ//G9i1Qwlp1Q8XahUbu1eRaDSrm4P
KmTZusM7/ffhVNQBMOnFqucpQIpimnEkT92bhgZ+1HhxWElAfGySe0dwaYoOlKPpFaVKM8J5zufR
nal0dOMhEDIYsIwPnOcbblXzwalOdaeJ+bWx6Uve5HCkY1LOFf0qP1TsJRHedmX9uk5iJ0TVoL9Q
dhm5SwDnFfz5Ax2+/J3F/SrgA7w23s/OAWx6wlIzlzxiPqW7QImXnHOAhMPeBPR0RNgQbwzCHfHf
/a2np8n7ocQRrueYt7lIbjtACqWfqXNonYeXMhgBGRUnAdRPYvsJ+1DYTuEkNJliCB3VwTEuePK1
Vxuq8JbnITZ8H+5WsGo0/mnE1TDzSw9zm20aFyBHcBAERqtUme125pSSIHmot/Okd8nDGV3PT+uv
qKFwKssYdTN0Uk+01OwUlXtw3/gzZeZPkhCBdmJp3YCoQtjiqubg8MauVpw2SCaK0aqr5SDOxytE
p5byVgKypdrWUTRq3rNWbq3D1l5ztpBEtas8mQGKynQhtLJ8RC1pkqb15T8tbdLNmm/TNZH85MYO
hm3kv0Jq8AISbcgP7LhZJ3OjPyhklSpVu6H1TNkraiEfdQb5v1DkYAxcWUO0mWZFUNnfSJgzV54O
Ps4WP0FCjiNjDq8QVzVF8gBKVcRN21nK3Rsv97iypXZ1T7JaM8quaJZYJSD8NziD5nf6aK+R/sYy
v5FECCUpeldLRUBpZIgf9bKLl2BBpmd8YJ9n5Nyax59ccsuuhhXtnGg8an5JDfc6Zx5ZyDn/Dfip
XimPvw1E3pD+tulGMtDZN/CusiNzt7bXCtThYws88KZORw93heIWFw0m0vZob9Ij76h/3mfhUSbw
/PhAU2LarR7Brpg80MmaxC7hyIps8OLpPFJopP19rlwxvrt5ArXgDxMUBX2QBtHGBmVibA9sHHRj
LBfshqDW1MLKJbvVRDiKmZxBPWXvyLmgCF8mR2mIMLnqjoZ11ol/w8kZxcVhNJ5MncE0lYiQ1XyN
ziQp1QBfk1tutJCp0pW1nvj74Ic6aeBMuHTwHb5QLxEdg7H9ETvooXzU3u3Ib4Lbz1iOM/dcx7M1
RRD8FhO4SMsup4Feb9VNsBDW3kJ3Oa5BQhxITIeY0ZmuFcqEVccsUAaXWdz2xhGA3/CiBI6uRCB9
tIndblsoJLqFCjxIi9w8r6nbqvPQnCExhO4x9vqxrOydw1ljwh7YkotZsWLuOOd0ICheO+mkVRIR
UzFhFRYmDSiHcgMocScdHJQ2nES3n86/lnny1gC1Kzg8OVWmDL+cifF6icWPTGdFqHwBQ0C+4gT2
S0M4PUDDHsnHWK2x7ymgQt4wcqIyw+L1ddjokUmqBVZng6s1kqpG/O+SpXdgyH0S8IWEcV//5UVB
tz/IHQp+pkZ881zsbVxxc34Ej0Jy+kIph1bcSA33NqDpnZCoORvZecAmCM0M4F73HqIks55TjaAz
rjxfLqICh2kjqZ/fteW2Tm6CUKSCg1hIJP7xB9i3fPccBDvkvbtrFkHsVRAhrakHcqENVmZP3SJh
6VtayBAe2Zk3wjs64sEmG2Uaw5HrkdkBznOtoChWKOPJW6ZqqlZoXEbJPc45mLrA0ynpsXrQdW3H
EGn3OP+rLIogJkxT5WfHdg1ricYDJ3HzcQn7MLLH5gMnErrDHcAlTod8Bygo/t02WTq5KGf95VUr
SsuMMdt2UeWElaVffMZEvVpEpn2GrXP7agnUip+xXR2skRSobEgum8b5A+xmgPXDrVsIkf58tOl0
B5c+aOPLtBiaNpfWXdETqwdZQH9zAekAM3P142+ulxaF5UO/MTLW1JWv0MDHZ8tB4D1El7lmk1ei
UxdMqoINQpNL5w64sObq4sJTmoYUjeGDU9YvQ/+QJiZjxZkWb6W9scLsvKrlfk1CFfdApQsLtJMi
HlKIcTF1JgDHET1E+GHBZUR6a+B4CJvE7HDzl+7qYn/mSaX6HXNPeGOMo379p55BVKCPiHLTYO0j
J0OHSl5z5PWRtRT2eOiFE8AZnBEL3ocW5NE6tAwMMHSXkXNCBGZgkyJTmMreDs1MYmdzYLX/FCZa
iddJmsrtCGi+fI1VP4WqSnBTLLWlhRWda4TSPy0Q6T559omImz4yiDNZYjLsM3Xsw/od6BX+87Nr
eyxbMuyNlyabxi+q9i+09FK3zeuS0t1edtmQTiGRxYEChBvFy1v35+PTgVkCpIaBd7SA9GAddy9u
YvY80zo0FadPNe7k4XJvbqc9puXZV1mpw5qe166xjq8bLaGhjhkhwEiMFPW2Uj5OEbtuu+tTQHUF
RTaiRZQjfInE3mmkdYhN4M2sZU8EJbb12iRsN60OjVTtk0KHqdFbyi9rrub0kuiVu8JBIYaJbYMC
JX8EyyBSDLl/n408jdYTvxRa71/PAb5x3SznYk62B2YjbTZ4AEjptbENeXr3oOdzP0tvVAlYwl9x
ElfMgi1A3Qs9Ox6MmATdT4edIQv3rs5yRegVACTaCsK4uWH6QyMsQQvMcNRx6+dRH4Dwary9Y9vr
0Uwz0FjSVCxDzw9pE2JUHZqhfr9ZJlLtkdmQjQNgm0LHEYj/zZ2pxI70GwjjamzOjuQI7AzU1C91
M4q3AXy6dAmtnITugLf39A1NDCF7iJ3Q8DTR+H8mkvTodC+lh8l4L4VS7DEdJqyBtytZuQkJRvtn
uaNL0KhK2YSjB9KMqJmRcmq0hbA2TBXytL0Gr63EVRQCgZTOvzBjHUbMq+NAijj/CB8Ci0bwlwOJ
2LfT7Kvb0YsKlYIB7LXI1oPMUgXeo9lIvOXKVnmdKUvcWxINjW4mDZvXkIsq1MkgJ6X0Vnggkshu
i39lSHX3asGrDIau/qlQiipZ8MfeZBPtH8HXO2BqiQfXGqx/Bj4Q7qe9ugy5PdEjihJvo6JSXGWz
lUopzHLcYMtyF5VskJ4170Dp7BGlkfCiIv8b89TyD3kphoVTvbhSoKVct1UxedBtbV89dq/UWRYL
aXhpc/QpCF1Suwg1dHcPHMsi5XIGVBmexav9brBifkKv+GKOtTnwa9lS0bpGtMNu3A87DHs7PF2J
Kmh5G0r9YMriuh33cWRNaC43vouZgE/Ilv0JYMaEQoVzIV/D8oK4O+bqoQ0j1PZRVgWPR9pG8fly
7+UUfgpEF/wlwwYemSJThNOveQ2a0ohC4nSOPl4tJbKm+/fO63ROCDkPiOSJFt8lGTl2mrtpXA3M
9AnwRC8zH2D/PwEy2FufW1hD3Erqm3vsgwYIA+5uu0LMz8DFrhC6D8B03YTLZ6iYfC1ADcFxzZ2z
NzNGui60gxE3xCqJmjBE8oFvpT+5MoYJN7bkbyvTsMavA6ynq40BqRPncDSeJCXkIXgWfe8iHhg5
GymDHybz1DByF8+sVepahWWaDoPeYLz/peCVT2ALMZIufhJbRkzz7QqaW7htQMiTlO5f3kwiRMw+
s4FE+OCktUGy799BxzGg0bogalnl0JngyjhLzTWRZJmm43e51guADzWY8D9FCzZSqS8FrLfAUNn3
KqLm0lFHFUDhFA8RMVzqFCj5RhvhMBf0HIWXrddzccknRYKeh39uGyBxtAeOWSo+P796kJqnWNcl
5MOo6mL5Sw8m7aQmWPxCWvpW7MbasiY0e3ZOlL5bQeaxTm0mZKG/4KH1KCX6Iq8e5NsCiDOVxAvf
CL/kG2U0Sf5Xr2a+U7T36SR/J8TRASY5CLUM5a3gurK69oBBTUf3bGA5rBadQoJGQAtPciU37e+O
zkYnfc/R2VGFGo6cpBaUXC7SoQzMo3cXf3W3IOR9gd1gekPfRutzzZuf0m8Kvs5o3cYNAfHfQD15
qZWBXtHO2Oyo+lwp5ZzfZSYOT+T/4vnDN4epZhT2D4Iu2Bvg/9NRNQ9bqyMxCeNoJ9uo1fmtcS1z
Gc6GGvTlAfq0r396jMACkXFTSrrXdRdB4j4rStQtylHBKWbMKPXxSSmwr9UhKmie0G7vo2tOMumw
pUIKH3LOu7DZwplCKnDJF7YQr8FoXyQabpGEibVZxeM1u87U7skZjCMXZ1oXqG+p4og5cqAjWXhe
I8JG2Xef1TQL1V8xxF8eOtjAJUqbJ+W7GWrNkLyGWMDHnvR51tcsSzP8zWXPN/I/erVgLDIweA1G
ZgmKarpY4d9BI5N735oWYteWipbupWtwxqszn7bmdyBQz7oV+AXZcbE0lojslJo5I8UQY9fYJtbd
DflAK3oL6xVN0d0FC3hxskS/pDyAdZpvHKohrQjxpfCB9O0LX18zU0BELOMYPT7ynW1O8mUIDPNo
6Ggh3cX+Jr59Dl6g5desAvqThEY/p19xmn8oG5bP9YYsF5Cy98LVtzQfxRZTJqfOT48oRX/KHuQQ
pHuyHQ2nazAvXdFp50NJsRmzSkh1ov3A6KgpoMkPwiCASiIlR7fTs9N/FRIVrWrkoW325aThP405
qJrYUm++tFe4tlb7iLGODinkyfxw4PAGY7DmL0tXAbJWPlpZjVE/PL5e7tV5A1LuETp7ei/Av6Qc
QA/d8PXOT7C5b+zBAq6F041X7kvKYpnlJsTzhr6ypJ6j91aW2hr1sTuViDpss0VCVO79gDJcqXK4
fleJ4s+dsTBX9/w3uCxMfkyCdf/s4+rN2OTqkIN5c16fM/tHSZwd/IH1q0rwjBvcZ1fcEyd2YnR8
TlJK9W2oVyr9hMB+dgi1sGTQ0UdOfq0U5ZLYbvGQxxP/Wd5KpBbhdd7C1qWE1ru9qjfysiRTcZPq
sKtrL1n7gQrSr4GnAPK2CsfUPAOHtNkTSsbRNMUPxaXcl1M31TvVs+nTRtS6EGBBrDWpNYDG5zgj
UW0eNHqTs3bewVVvgF2VjNOM5M+Jcia32Yh4tPhxEpZUN09S5rTxzaNHYtVIHcN/J697Nnj8YnJQ
0/f14wPQkYs2a02NxYwtj41HdzsfCZ0lEQhb42dBnxmGLRFBLFv4AFT+zPdZd3Jy3z/DaKYtMg+q
ESwbfFaZIsEGbkcZrsOw9AWAd3cmHHHUlSGXYN4/dsk27XWcT5wrcUbRpc0S48a/350/zDB/7IH0
TxFIOX/5X7zy3EHuL1De07NxxfRNncfdYDF6uVasigc/sINHRI5fIN6dpvpozbQLgfa2UlO7bdRD
EqELIOLRBGYDHMvmFWkO9OzXQfGcrgtTx6x3feZIk1RJp2+0BymxFzBLGqVS3HrDk4K4dzT61exn
qIkOOWXTTdBhd9kSBbnL7Dtn6Ne9dDYnMNwaCVSqO1KBUaMs1V6DySIc6xkhRdzVeU0q7nY2OWfL
mYfWbNeIjzFQxh/5IKh52+339Fil6A42lDdBp1cHooohRyLSiXJgpi20ifptFJcDW34kCgOFDhBE
HccbOqBRkoqFets5OW3xnD9njyoEQYqs3+VHvdbu9nqWX+/b8kxbJLXFNBJxTVTQI6rBchpMzAQ1
VgDPtyG/Wk2N2gO58BYNYT36Y1PeB1S9dOltBIqL6My4CBza0gqIi+KjEwYILoyr4bciriBs9MOE
cbxQcYPrpmGlDpuoEKIWVavn/uU7owK7dNoOkGfvgQ0/QkCR/CT+iVd39T/mZXlxNfD281g75CyF
Mx/S8qlnDx0ZDWZU/73srLFuJwO1ynXPkJBvlFf4syarP3I+WZm0pTpRacc+wXhfyDWJXI+bWxKz
ABPR1W1y1tD5NoRY2JaiusTTiTk4ElA+f8wfHf/DTEYdpUmpy+cHkKH5kb6ClDbsZJm5HFmpLTq0
QPrVEKnPUkpwiKv9SKQ4LPTQWEAz3ZnDXP8or7NJh7uW2XQ8w2HstxQbV4QmrxdtzNA6zhDaGkO4
GCtZZqByQEEkVbNvBV8dJlkBMe0kyKYF8ycgqq3b7+J/1YjFxKz23RSYO3CZv9UtiYfc8LpIcTvY
JE3rzVsh378OHdSF1G9cpu+3FhUyYJdmPD1MgVQNrp8Hcg3qs12+7TH3aCAldSNC0nPOHdpp+q8m
7cMfXVbJ/j+WY7X5KLtUrP8PGyfBNnHCTPJYhgpd3YA/HMc0gZcjgiT59o0SxxtLNX3kUDfPKiyo
WKwWgeE7EW/WIMP2vPAOs3qKODMWj3A7SHcgkr1u+q8b+plz/yUEfNKTGdtuhjDzlOKvgDpBe9kW
/FXg567Q8Gsm1dX/7yaXB8IpfVqpS7uuYLmmmkizLioc7tL0TlcGHM229aN3vNrUGWfyh0WWndz5
jz2G0/3UyqmUTd6lBILeE9nAZvL8a5UZ2w0HdF2XLe85vbrA++e+az5InZGOH2J4dUxl0i7VmR72
UcV6AbgWWC9NrmXL+c36Dpo3PG3mr4nVr308oTUtHl1VYEChcEshQhGulOTFHPFBYK9ddyWajSzw
LTuvT116LwTm/4sOG9HDKxUXn62ZXhr1sA54DarTpd5dKeAuZTJ0/93UzCrbCwGrZVBb6pXdQ+Yf
IQwqjbyqjYf/ncTweiunxtuN1NYD+SLNaUAuPZ8elMZqUFPdb3ODTKNbOd8Fzm128/xyUcZzeH6x
LwQLXTpWabbFRpKnI/AHEfoIo0t6DAdE0gjDlykyFB/NOaAaX/BJrBuzx0WUdRSLyTdpMNmLwX8c
wfWviI2+bxpvAL2P3zuZBp5xsyIJGoFiw7SAZjwEDPhq9c9k2H+Cgv45cZtQM6+LUsRbuIMpTU+t
N+Tc/idZPlr6ZLyCxEEEGlWoWTLjzRi2lZygJ056bGDK9xJEFvqshKU06XORlEcZDfTvL0Y2rdSM
zbOhf3OGIdA6dtFI0uldFNn0LVpFCQgqDFJFv+1GeD++V70TPMROvl6AKMorIWeefc1rAJojUtf0
64lc7Qbktd7sRDJYKnCD/xiOV31jXfmFjSHyhZTtXvPDY/6VkRPjHTT5ipZNBqLnRtZRzP3ZfnE5
4LjAkYylVm2b1l/IU6SYbx9ll0FOMv2mvZs8neohQhnOuFO15dT+dfacPROGjPq9r6Feg02NpR21
kQrXscn08Wcdw4u6roMEbh+VCUNcboR+5Cke7IrHEs87KIQLVd0RBhx3EgpdXmsmaApGWMXlS9rd
au3gMTh+YTBGQ/45nn8PC6DgL3fRZMVFaJ1+bHqRJTTWJFjQHHtQ3btxgTyt7xuTf6wmN1bJKvuc
Tf/q7AG2B2JIERiVsD2fpZs2iNt8QcTxp6l30WQnCivqrdtovze38x3AWB7qc6OxYekv0D+8Vr/y
vuZPpOZApjXhoidqfboTWp2P2MHphXt/7HLXINStQpC6r+asqUwDDNZs4BkI8Q3jW9c5Kn/c5MlV
SnzBc01oqz1fhI6LcFesdxByhcsYPGRa4TxW5rpISQzy7SWBmNn9/DeL8gHOE/cf8+CU+0Hh/Ang
ZzMZ9/TXG3lqaVq8gtC/FzEHem1LN9J2ALc+WO8Dp+SMi44h7vWN7yl7CIFbrFSsORBYGQoGhT5w
+Sw9w0hkNzIwbrGyXJI6wWVp1+cFo/aqTn9iW2vOPU1gBHs7+JVoo2LecgOydD74Z2KtcMQwFGbR
os6C7Zkee3hf9YuZrnJDqcxbZmi2goO5Olc2sK5wfleXqAktKyyf6H4jiBxUQsA2aNjt2yMlNZgW
rY6tqHwetGzFqaRUjnP2olnIXp05aBA7/hyzRduXIc6udBOnMh1AnMZBqb/Z7FYK6+lKENdnrLI3
JI+6rV6OurSLBPRGZgI9gBAgZr1Dx6PHKV3vx2bqTtB4GiId5fI2LQ//IzZKG+B0LVyK/7ZoZK0z
kc6C5KHcCd2rhpSkAyLMsW8ulzuAN1F0X2sflnL4ScSiOgeBbgUJrLMfZolaZCiHB7+66VBP+zya
BMigYeyM5S68VpTnFi91n82JVIapi+q+7+5h2JvLYlllSIrpiFxxbBIV0ltohpupPe8V6yLSN5xX
81AHKqb9qgRprtrANLEuNfwmpO98MiC8zi+KDNkV+RSrhPnwWw+RAHleMXNoLcSr5ovq5KCT1NHo
NllRpi77dIGzfAgBl9qcHSRvOlYWNuxjb/u5/X3OWdIavZFml0J02DvMEYR/aROXiDLxiFHJnVB6
WV0d8DavCvgGnphkzeHZXLU8Ow8SJWAU3qFz/26HX7kFfvCDPTbHzydlAzIu8CcBDi2YZiR8CHs6
ORE0g1qylLbVUAFp5BDSI2h/oi/CrnLP1XAJENEF5MQZJHvizg1sWSyVAA/K7JzH+7Ohj+1hV/e+
HvFaDrkWxtA/B0Bxa1JInLP1r3U4gbD6/pOONXdS7OUK0wY51BLaQR1YqugTv862bzf7mzreJY5B
ULdCZG8hTOnwk9gx6SOC0MV9rFkDYAvvHXNRxWtmk9aby36IThzMX0QB1CG6z7zcgMXualMK+3Q+
JPccPbvymmm/HPfUHitFYcGhppqigdV8nPTYKFoTcYf/uMVGkM/6DD7KVqWZ8sX5eqLi2FcaxeB1
lzhb9Oa6rsZSUrf1oCq0ErF03T6pCEfLF0h65hItsesZcI4GL4TVz/D1BzQnAA3Kt6rZ8tpM8/89
MNEP9peGsLAf5oKCl4d/H2pvapp/tCEG5WAlw+W2uzzGjqoYWIqYaBrGhkt1aasH2L67Jaat6pKE
krLKj4YITNd49bgfprXzfEpSaIb7o4f1JM01PUI5kHck+xHdNbOaAULkTGG4QEkPLom6QO2Y0a+1
iTED04hyHpYm0hEWnKSmvDosuQqB9tdKB/JfXhSZeouKrv3DLXvYtQu9gpeO2ahPZ/K4SRKK4u9t
9Qfh448PrOSh0++84wL975nSWcQ8TyKDqQPdf+2XBlou2l7AjCfFX0b4uISIAx9+ThW/uQuAMcbP
Bd9ZoJMwF+zlW/mQTcgM7uv+ge892eUC2HYSQDVGgLP324atBnhai8oK6CaQngUrQkko8OfZOkV0
HsX8fh+UIe9yfdmBOo4QcPD1AWkmJYAr9QrlzmnGQBjvkclOF5W8WkTd2avANQHPeVzXQKAACpPL
2andf/U16EnZuJuw3Q2Wu8d9x3CQOdOYLNiarkTlg4JqEsngUydBgewFLczYdBvEuzmdvKGUL9ig
5IL93amVZBrwapuGyDbyBjq6vpQl6bbiqbw0l0/eVyxaAlgu3LOlofnrqeU31hBBDK7E2h+6Ir1T
6VMuTLNzILhjdZxD0gRsZZWDBUP4Quf8EjSUAK3Xx6z0+GDdupsigQCI2v+MX9nnIqJzElG+9s3X
TN8sVkKn6J8Pg9n4sj03IxcU3HHEXvCc5RTrgEVsvM0KI8AlHhB80PABZyQGUjQ8oZShWqff5eQO
wYB7pb4PhCNFYyLh9/IEuVpm++THClrKKWgfNELrK2fig7FStNt4xnfbgetn/lwreFG9oUbATqL1
ankyFkhZzgq/S1VjKtMsoWs+0p7f/LiBza6PhYWf9N1JVOdXEfE0qm9vwBDoDO56ncHt0+JRSrHo
COh3nG6NXnLbKwmWdSvNnunCGyWQ14LfkW31jiUccUqSZCUtl6HPoxripmvgSnLPAU6jj7LoCPMm
qvpa1uwE3+d5M+LZNs9lsHtX24OzUcGIe3zxPAOQtuV/5vCYO6D0g/jhTorpiTNIk45Ljs0lnv8N
+/+cny/PikvZgfn/LIE6QVVfr+dy9UfVSkvdHmnEO83e8A2yXLKQYOSLhH6AGweVksieb8PXQS8e
/zLXRbFSE87ZILVAFGtnO5Q8KV8uFiBkPwMpIGhiKk4ZLcUkCD+QoqVdVcXs2UR0uEnPIfDcLNGQ
dJfxWwbyh1JAT0t6DlOl/eZvrY5FtVY/1fiIEMSEtFFY/Xuf6ImAoUwGQG+i2wKU7tKHXxgboSpn
hk6//ld+hyd+8Y3VHcQkBTNSzdU6Rfbj+SmwobOJZOoxxznwS8B/3vQYcNAQzER/Tm4PvUxGV1BF
ZwZavqIuEYEG9ZK3jXgdAHs3wBNip3N2Y/6ZiOMSCPnWRpD85HrtupByxJ/ou8kfgjBLWm+vFBLL
tZvT5TwfHBNgdRrAMgs3+oVG7H1ZjD2W9Mm8SOZEdGwm8NMiAImQB6vuBjs1riHSsOtWJUCfcGsx
K/6Eexhsc9ICcYSV8DKEYrslR8Ek+f235LJzxjs3YJKroKYQSpET9y7pZz0bK3sIvJM8re77xo4Y
WNNKAR1fLXTl39KXqC2RHqPdZB6xMSiPzQHx0siKC1aStOdVFmgzeHdC1XQ47yoPVALFshNGQAAz
ZqlO+zkTH6pY/PfrX/kI9Gim00ENq6ae4HJpwY81MN44oTJY3guWlO+exaAxoxJkaY2NdE1aRVft
jJf9bHPY3MRYAD59r4h+z511hI9LNx7sB/orCP24UHAVnRkV0i1man95xL6HBxz6ipZ+cQzoNe46
zavz+sHrsR+jCvgaxETmcRaVLZ1ZIOl8Pltlju/ce/T8lFxJOlfQ2DywCt+AefMOViWWCF56TnG8
wINWSMzjrBmxyjTdvWBhPSBnqa7TgA7/od+h5xWlYxx/q0RRQzDQUJwG3kjqEfabGC9I86JkCaNz
4EqlR2df/18A0SdG7S0QsyhlK2EWUVCmKm1sNqvklVntHminNwDgiXh+PevC28d90wrlpsSkkYBn
vB1aDihvb354nU8OIUZJ/9r9eDaqdQlCIkTBXk8wkTVKjB3H38g/MnyH9PO7RCDJ9JbW7sxk6ObG
ApMVFXoQcGynr+BvuSM83ZpGwOwnzeLIhAVw+tAQXlMUmHuONsIY1PZsuvF/yps6NzNsqDZbZUA/
OB9Ji/4QAgX4BMO6lFn6/+wikEvMeq7HJwsJOcDFQoDzCCoeX4hzvS7J952tT0cyqoGNzb7srNjr
MWXh4dO+aUF2snvYyP/TngEC+RA/ROjDP/e+4jAUO8exoo9Q3ERwBUutAzZvgRKCNf1IkhD01bAf
4OvQTfp1mUXJLeDF8WYmzwLF0dCno+BUl8Dk9w9RupdmQFv7VH6lnLWu0DwgG3KO8PTJLC/sytzm
7nG+AaEmh+aYxyHeCMArKM9K/w7UR4aTXYIAq/ZnjI55Z/DYKCnpAyfORD5vqFFoihK7O/KchSuK
A9ixMLoK3BlH4o+c7jN+naoTHSrUTDDjJVFJB9Opg8iBM7KlOqe/o041iUYoB/5VCmRI0Az2HdNB
WzZcIFV/afnk7wo8jMsxfLgxJkHgGkz+BliWb9iAw71naiz4sJaWBbafJn5Vr+6Mm0yjEPwkMExU
GhjlCDu6f2EntQH/eh0TziTTN27DUF8NPOzBALG9UYr+XlTr+phnXXE7d67tROVQtIbIgkqz1hgU
cEVo2dJ55ajg3OVtkC9nTELSVngt5rfoGcdcz3wiIaccWrg1OxVoqoWIVDCTbeyvMfVJ2ouJqKxo
ErXJFh05RCVn/7GXhcXKjP/rq+hw5gQkKcDsnQUXM25RtxRvlmSI+LNQedHSCcTlMhxE4mJqAehe
dtruuNQUVXSh0AR+LLXn3EA7kA/okPgWKON1klrnz8nAPXkjnZz4fRM67HDrzG/d/69gZfRkRiMU
dMs9JyJaH7ELlvO0q7BR96LCxIpozbJbWo3jiA4+nq5tJEc8/Qvs2AVzLuAzwFlV1hj9pxwJNfVV
DgmOlzjoeHT0LNfh8yBy/Qo3i1CTpoeRkSvYAr9Wvv5sQXjgMBSGyoCpAxVzVozYHB9Xpq7kA1Lf
X36VBFTiyurgsAizxcM4HsMfno7bNGTonqB8Y+AkO9w2dZMsWU/VYQDIQKAGI5zUkbdhuQw2gtBz
slepSMN1fXLL4KkPvMOqPYvaFN6k7+bRMHSRNuxWR9uQJz+3rj5ZS8CT995j2FJhjk86fi0HL6aj
icVwsWW/13r49BpSxV7a/9xzSXXaTO8RCSImxJCL6x+xojoRzcsrRGHh7G4vOTXfjGxXBofUGMHJ
gn68TTseHyBtm7JskcCo6GjhERV9IlRqKSfetDeG4bkHMrQWAVMXVWmK/6jtptJXBVFuhK3IqX9+
f573L43285UsCoZQva6EAFDd3zegFoZyjkctCsScLm4EW5NoCYsDIYeuI9WQWPlrxg7FeHybZSpA
3W8V/e1VnwLTk6ZY+FEsg5YGctJOJdPG/hgDoNAE2qaV2dcNBjtaxmmwOykVqBmLKh5zbODrsGcF
NqqY4RXMy+lETpY/JX1aTjlvElIhv/9SqDp7u6/fFVBCEFOgva8EYbuEzFkag/bPaMEq5Z2sLMDH
1wJBK7tQ+X4Zg/GAHvAQCIkTWv9eFZFOY5Tup5mVVDnJIAqvh+KqGE8T7x4iYy+gOmNHsfic00m6
vEghRC8LCVTyNbxobGnTuzz2W8GUP2lcfJa0o+UEpSX9ejWk8GPGhUQAHkfmRPJiamiIQ9dKthQV
lTCt2R4dkdI5ja43Noj72oHNI50gHiFFZ3lK4ht1nzM1QlxAmet+O4hVxk2v/Jr1ddyFm48e2zQg
HwZBkKeyxDU8ETUSId69PRNJejEUE4UbC5/t2PbByS43HCSTipl5q82IiaqR+pCbdUPAtHamkSC5
Djf0/mfbEJDcUCc+Ssbtvbjj5kaZ3u4Y3pee947iGQbfHZ1Ed9Ngnx3QYZG6xdbmucAzGjqR1o7R
y8HZZ9HxIVpfuSLaPAbq3BNvFJ3t5SCOYA/lh2bT6ilJlPdI3JwS6NFPa9BkhfsUwtIZV2BaCadY
2BQ3UBAYOsewa9BxK0v8D0cR9hJEpN9BZ8/cY/Ywzomx8Vip4+myYwEywmXjnHAoFk+g/7FoKI2z
W/IY5KmFosN1cngvMStQwoN3Bp+6meg4bINfjWz9jKAHdlPRtgApYnh5uCCb9qiKxJUGlq3nmWiW
X1ewDeqbp8AZvRLcw5+aIlbsT44VP+Wl1y6Jn3be6YYcAQDxPFwaawrTS+AgKy6OdvL2JwfIZG0f
KhRF41m+tPkaIrhuNnvzmIIYzSPTxoaehzgzRRtvbwpbkIUy4uguVXi18cPT2Us9+P7LPzfoSHUX
UBe0N2/o8mGbVzLHz0uf133LXXtba3u8XRFohSGCR53XHboMboYxPtBEJcdVxKax0PMMA6aXlikf
uGZU8NXxdHz/3+JBA0/IQfS2M3wGnK19jvAJzCyMBJIk14zWpQs6apVX91tmdvtdevyy9wkpABfo
r3Sdb3ZXFbVtXwKKRcP39pC5UrSplsqAOBEfh9+iKPaB1BjnLhmbNUBA8O1+nd+4nvl1NyARDHU1
AVq7xT/T1vvRdqgO0lF93bO7rwk0UVi4s7CBDSttUrUPQzlKbG9j4nq1UDthIVaNzLxq3mzcLRmX
ZXXVxl+zsrEFFw48IIWEZSktiDGff9E4ZyOMfNeLYOFT5FVC8Sh4B1W4wIvTOA7p+VQdxSmAdEpA
VxYxmvDepRKpyaYOUpyBXFwjRdMA2/CXuPRnIydgayorW08x6hrNkCd5CK2AgQGG4cU4oivqN0Xy
L+qts/gZiX8JfKpfFTSDR6oRIlpzQIds44RW0UgPUt6zwYby7r37fx392ICpue8kkb3UxBHQ0XF2
aOKUfxx/EqGWwy78dSLQ7TUZjbbuxrNYyra1LYLm/p+UqwAmShq6wZLzKOPDIUCdy/BQQ46rZJQ0
QCMogLyZywJtZ7KF2hyavGGXJ1rQoxqU61KOrB7P5wYe1AJTnAwobUN+0h5t6CEmKcJxjju/iW6+
eJOGVisolJ8A5/C7DihREq8TKuCfxiD94EMpV6n/Id0SeRlUEgfVjHLfAypnba/qpQrIVZOSp/TK
uqrDTls9Y0VA5GlyEks5XgV6Y425HbmhTaJ8HyWPdsBCIBOKGyAjqYn4ZGIhsVK2R3sanf7jrqUZ
ilo0wVdV06yfs33E7B8CmjXYVN1gVSNuMyz3M87g7TktBAxqylDhMV5g4fT7LewSRcZzd/5f4bFA
/3Rl6sT71WMJ9nCkWzhDYtGmPlaDS7k/PVLwZdJUhCAvtskBRQJEwBBnZ6FRarJmn9lLNZosR12C
3sUGsWu92hr1hKiyQit9AU6che0zJQh/YjzD1yq7m3n9bCA19lwgwKeEhBIiTfWVxJFSRNNiKrcK
Ek398XzjOPW654cA2ervwfVLkVwfSp71zNqn7TZ4k50w+pok/bfFc9Bb7hvGHe3UPIFq8UnE/Iyh
tjVG+OFxOjXIO3Zbt89WZCV47V5aapesHdljORhcY1IXIp5uWGhz3JV/9t4i4z3amHMrSrZINUTE
fduUGh34ViLR0ADZRRI3kxsOjLPOG43YvkpbiYI0Q2H36uauoo3/tQVlV5iBBiCVmGoB/VnWQFat
4W74XKnz/7AWygPVQwUdblq9RloywAQ5hb5jEnMr3FUcf/v78LwY4l8RYMqN01TitU8ZQswQbz1x
CQmSOWdF8NQMKcPkoyPPcj96ATAOkQyOnXR9b07GLXDySK25DyWKNCYN+GLF7deWDU2hb0dRQ9NT
bOz3UDsUTlgcSmdO90W9zBR3BolRcD94PEGRAUwq3DIvPA9URPHIvJQM1R++G09U3aVran0I5amx
V9yXvrGwsoQAA/q5sH5+LoER94DTXwgMEjVffBvezdlcFeLKBBFXcqLu6T/PgwV+At9hK5BdfJar
xa8PkaN2lREkzq9iQKG5VstDEDfHxUN4KYuOrP+gkpyYamSlVPFzpEJgcgWnwoOrS8S1q2QHWCRv
PENeZk37Y7rVZaj2E5c/0dgO0uKpsRE8rJM27bVEzaLw6ldm4AWW42WeoOCtwsex5ztIYBhnfUcH
qkhuhD1ymz314b3OT6TnG9/lI3DCynAQsCEJKFyb9o75VjpMkbqNz1j1IRyAtkOjwupkp6+ryR/V
KTrNCoR3uednPnoDz85Nq41ri2iL7h7nOyq4n6h2Wq3WrZ6C0pob2HeDlxGcQbDfRk1l6imjgFwP
smmM8k5Xs41kWj9Lhg3+NFDsN86N/TU1EdNKPP4CQ9YlNizwo1pxDmSfqxcw6hSvXt0zfa2UAEk9
TnXU3Zl+6ksdgaE5H0Dkjz8dxf7Znj+V46l+hkkNutxj/Zz0WcjfL1ASq20S93LO4V2g4Jh/GCk+
s3ce0vOJrx1hYAWL+3s4hJVo3b4RRD3HSOoy3AEupD1QFyaPB++uWwXJTnTBfBWSSLxYJDS/zm2R
jYPsQnV0jfwER4Sez60Ow4rOJswHCRFQdbTwAEbru2WaURQ6bkLhGxm2XPKSbm/oEhpUAw1EgNcr
HuRhIs2qbf/os0B5RD1Ro3WuYdBVgEBqDPYwfuUdLsKEmp3aAAb5PqGCPqBSogFcleRZsVGX6miC
zjuVGkMYCvyFRy1g92kDZTkAWzRaV8z8tDfziQZf6gO2GEZekBeMcfzivZPN1YCCenhxz3FxthTz
K3MNonxrBRX0TdTpnkQcfjnGHkOK8sEZJV62BwIfaPhh6r//R5oyYCFpumTQTDm3dnSYVhOc4m5g
Rb+rUXJS7UIPUgbRWV/ZZvYVJDuUx/Cmfwn1yKNGo7h+i9D/uAqJ37SwKAvk31WhxO/mTzQ4kc2N
/Olz24Dq5ku+AXms6DeD+yDHxChzoGzB256iBl76WVR+eQQENAxh0LQJp0Kv4ifR7nYpTY/uEtRV
wEYykRjbyGPPFhPEFRch+CXJuVKK2Te1JKGd4e4l5enlT3VPeGJHJ+u6pJtctOwmLOMvtVBsUSdz
HPBYmG1fjQHJhwwFPrLscEWEqCKeQCkakt4QuoToa74d5wEMNTRrrcAzwXyDIXEzl/95YOXo1szq
2WxvyX+q8/eBth8xQCjV8EAx6cMGjU7Au1+Hq262hIqtBYyDYhi95ddtV2l13qMvadpsrSjBAux8
IJESVetNLPvVzqV9YdEZ3+J1k6e9PNQqiVC7CDEcR2OWHQvZ6vDsfBBMrtC8c367PwTiSZzDEj1C
nT2QVZIG0UC8RBYwuIK5GcyrvSPSchDjPWK0E7fzuRYjaFFTF6kjPuo65e9lpElRXA8yyC59Uk13
BddFn8scHMofjnb4+IrkZvem/O/oppJCRm9J0jJ7enIE5n3bEVTAqhbHTSf11z+Au5nDv27NWtI5
8a6ULcCVKx3CAzagDiUdehHZHQTkBbZ9rya8zsz+JvN7L6Qbvxobxn+tWOPC4QNk84njglUidxnz
pXZGl09Na2sW9KCfZ3lh1VxkrkZPM5erR1gGTX0AeTCFWMcxG6blYIQMj1araEZ6xZOJBT0fu1YP
18UdghTUG2gi+rA2srFmOFhjA/f8ut3Uuiv/ya6Ra8S2ZyoLa+oSknVxDH6Blk0w1RKHtiX649pp
dGM9Oi5glzPpiUA0STCjIevKyKi2iP2XW58fnw3IF8K4JbCZPoYi5y/8eTgWusOThBGRk/GaEomC
CF8SVGvxJcSZbnlWwlFpr2YzNZBfZgkEw47fQbTH3tyGXi31ePH2JDrzoKd/qr9RNotQ74rs8cJg
8SLaY/jv3apgIKjYJnoBXR6aVQ+2qxQUVOV0N5yyTD4QKxETB9mkvKuX3PTttD0Hy/dW/JSU8zDs
EoDWu5CAvz8Supj41PPMElYC9uGApwzwqAV+Py4H+770ECmGde5Yfw92UUv7Xr/T104Ph2JVpFwK
4Mrn0ERgojTYHu4RY+08jrnN/+1hdN7+S5L0WxKGj7m+P3/i9JF/S3qgcntmzTGKOpNeOeHqsiFS
kyhJ95AY2wMWiBTynOIFEw0CJ2wK/vxv+zOoVnzTpzQ4NJ5b6w0ef284BlEH8eMlenHH3HVzAQTg
mlOhlPXVVdvZXlOz4aTW6G2yjSjfkjasGc9Ynm9fwcgDoOM/n7SbNKMXmXhT9py0V+1RTalmiit3
pxvsffruaPCsgoo4+3ekLTO1NVaKVU1nuS5njny5vF1lXUmA0I4X25u08ADq55eO3S0RCZENYEaR
iby+/EwEnsc1HFkHzNxF8HJrY4blP9RUGhzz2f0n7qbqckVPvfDwrCc4+rq4SFO0evbZ9k0yBHvD
LfFsF1o8rdKaxd0G7HLLR2D04GoUPY0tnCkci/a8btUm3JXzGMvNfFyTeUfC4Fs/9WF/U36sJATK
cH9oXsZoSMUQWPo6SpYykTNrVpBvqDbP+wI2jw1BAbsha8HfyA1ub7X/TfsDSyXc3w2ukVjaZR6x
b364Klfl/XdMzpYGb0fakoAAB0x/eP25LsnW+L/98+jvd5iC1P8gIyAWcoeI8JOGO9QGt+62JBIa
BpvHRxk7KG/NdQQDBQrmMXdFGA/Eia0yrdU1Yo7mXTV40qhvAHFtimvileFQnSAzOi4HX6l4WaPc
te0k+83vRct/Yy758rsq5Kgc33hZHrLpsYPV13f9nLoYzu8PFUaSU0pdURRuvbtcDpjgIUs/SsNc
B0ig3FFl/DhPNvy9uddeGOL/23tGeumKVKrzeS3ZHxlPV7btlPcU3aqQm+hMyV9IAfwYa+Uv+hVG
HQe7yTyMMwRlWrWwOo5DQsApfnxnvFpkKwz/CwZmokFhSw2Ok1VmJ+Kx0RzDO3fdlCBWLQcCijUA
CmsExlC+LZCwicFzPMdDkbnLJLUlI4e8uxCkREwYOfR2c0T5ihm4rqw6GA1RcBHL3mRx2/+LhKUu
eRk/+heb9yoyQkDEgfL+kyCmqiO+Te6SEjx6cdvJ/i532BavxjliDa8JxAmtyuqopkWEoSdiK1fo
4gc86Oh3QRwfm3qAh3hNU9ZME/I5E5MVvN+jbP4FY6QxBnKE8Y0bnYgu8C/RuxyZUDKItqP/a56E
BuL1iCsi2VOcFFBBbew9iHCujVCqKStVg9Chjyqa2EkxMSL0q94OxUgHKp/1ddX/YxwmDI5eN/gt
Vz6omBpOmvdPh7e5CFLNmwgUfhmOsoKot4Sm0t+XKGU0gedaNJcQdObdq0dFJuqMW/O/9odQg8az
VnGzLJQEn7Dizrdu/ayJgydTL4zbLx4o5mrY9U9Ow8TJUzFjG+155ru5FtKvKZQGs4WBDflhsygE
uXta2GqWZlTAsfs5KP2K6r6mfe7Yt9aAgYuTV42iDr9AGOEyRi0EswI0SC/e5sIEJQUgmOevOZWu
TsxGlA92IKccKQ1Sy8+/nqz097+4ijmkeRLZvttYzjSzFWzJ+glAIeLYbL4AAQu2/lQDmeQyE6dU
0NQkHBarPT++fCLqcrcnYhwmu3k5k39NyMGIW4XTy4JYcjRQHpMBWaUPh0kXPgK4tUXtPsvxHR7t
wILcW/EVLjHCaDpEL5fQ2/F/rS0TU17K4AXSfFqTxCEC0nkDsvQlXeQ9r/GJuK0weLqW2yK6HH0+
jGnmLFIrAzUEkWkmkRlLfjH2ZofMyYpJhDsYMYLQ5PhtX2d3drLs0xw08/99zUpG3TpYpAkCPRM7
Mjxq00cZz0XYPffSYK/jLISRoUx3O0/c+UXDlC1F1R7/Q5ODlip6PM0ECo5mnvry+8MX10rNE4y3
wdusEq/gE6XXNFjUGcJPR9LtDvzxx/aMixzYz6wQqFhnfhLf70j3xzwqTAXTvr5gywilbwmXv1eU
K8WlgQ9MYdEBKXEKT+1WTgI6zXwEtjx+LsG9dAdmvlKMBdE2Ru+cQ3JvL6OwW/KDWJSu5pYiZ6RB
jjCDG3a8PBlCvNF2yOSAXShYdcngn/HZ+xJluhMi7nOAvA2GGYP7UjirzwSFZgN5SywEn6Mvbtrn
zKycOn93GKNr48etq5riIj5uzH9lSwLOrYbNDPYS0EeGoPsqIsS8STL+37PP4SRADsUamHy5DJ6Y
voWhWNe+qZkTu7ST5V7K6gvWzSmAMKrH7xpvuChKNWsFsLahSYTsbqsS9DzH+eEmIuTA8TcOQJGb
/vE0RhuVIiBkz+qw/qzQVEtsT/ux2BKBbsS6P9rlpb3G/oduVPHoyRbfS0epU2x6LeV3T0/UkuTr
LHQ0ASIopjSHaCFQR+O7hgZI9V0RiILIIcZP77pi0K5Tzv1SV2z+gI8JWwMA9z/UoPVRvb0VGpnh
5l7KDrDWO7UNH2nJwvrVUcRlNfcHpDAfpMNxePNxKXNFJlCOJNhb+tQS4/09ZJwP0q+v6XCDb/As
bec1IesEH71aN7uLWSYaMhvW6bGQedQaqcO8pVqq1SNLcqWPV4qr8o8qcM592ySjDsrdU5K3ZWUu
qYDQvpB59bIkGrALCXarGaGyvKu07gj3PEA8aRlg/bnKtZSsG/y2wuBvAS3moaKLRhsUBy978MTn
e3x+M5Cmmg2f2+Up7mWthMRClUu73TlYP1GpF6TjandxhOJLwUQF/tAgSS74vSnaVTwac1g3HuIh
D9LrM3eME+iGs7+v4lFmZ3MKNWzfP+GqZlnvdqGbgIxWnGd00HwOFqTG4nPw6srVkZf43jiUAmur
T/v3JXK28rmKBp5Z2CmBvomCJJehe3l3v+7wxshIESyk+gCQXsd7D2D04eGzQN/dJ7ljeBB6cfyc
R90nNnQ3cWRE3Zfys7RCcKxzvrowJmWGcYf07zpl825MGshXzlT+mZ0xgKL+NMu4IXVL3qrYAd6v
WU5z4+fBX9LwuDFCJhJTTHS0HCh+1eUCKNhXCoCRYZU+xrYUoHzGQ706eiR21hLAIAOjpOHIs9ny
D/EGa0zXxYKuuAzGswoXgt4oQ6qrPBLgEzjsVVAGQcAoa1JQ1Zm85gEiYs6Kfi8cxzwz4OnrXBzi
PPzxXLuNJ3/0n5CIbSa66uC83aK5g9AIph/QwEm6ZEQ3ly1gEULLtlk9xFm14cHE8RMX1cOiDHdQ
+3FOZoyG9ais0qOnKv7EziRbgWSHgc0NVRYuJGdR6mRCe2+n7Rza+x7ew+uzM4/P3FQFI7J9F/Ov
WDAcGY2H2EdB/JKDdwLHsx6Qi9Z7NQCTEV4+aA1ipOnwK4pZ1/Aw72K65UIscklGNczOtvBwPcN9
6S1D+/EjgWTxUEbjMHMxZVmcoTJ1OCh8X5QWaKbY+8DUCyEfkuUdRvL+pHbPUCd6bowTytyz7l5o
zK1hqe4PjpWXV9KS1R86Slexg7jA7FVyJVzH57hMlpvO6JA8GZhAtY9BfG85RcXuVzn8LGTEJOJs
6Row11vKScof8hxGUck6KybkSr8ROjBz/c3yYd4i2EFGo1y0ijdEEScyNsRuB8OHRdaIbxZUambp
h3wakZwcfGHDLdXFNbYUDPjZu+sWDVDWjgZcxhkRLwRTmvYfHk6xJLFI/cyu6EHHEZaRAADBPBfw
lb0JnguEvc9E75XonUHG9tec2qCG+95hAAl7aEqXkdmhqYmA6OCp9NN+HxHQzIsZl9LmV/40VawU
aEiXLNW3rLDbgNy6rcwGfeJPANfRglWdwSHpypgF6CfF1Az82uUGN0rESeC8R6tlhx34IcpUT8C3
MABM7iFiMQSyYTUrZSAvekv5xyCKpYw+HpuIICeMl+7mc1cKhP+J2P78v1r4oyngMJXJVLIWfybn
z7QqvIUVkAfx9l18i0obw0268rjCynoX8aaj0kD9P/gqZPv4xk2Wz6jzB+YL3XzBUrptECUWoUOA
c6MIMNB9+vAqCf00CERsxPH99sg4y8EGiClsXdUijrTYwBJO6MAK2OMbPz/w8APGw0eM7LT1zMPk
wbRwNfNTRbA1HKAIbD8Wr5FKkITW/OyZolrNEGDSMZdiFw6ToBxTsnQxZdO98036aarInCg8t80Q
DwpkN0asMyi0c3tqiE+0/amUiSRBdA8IwHIyY4bOT0g8CtErUoh6AGiGOrCjCCnZ5Ltw0AOpZX3m
C93cWa+/UZU0OgYKSABWzU971HxdmQH97V8tTcOCDXj6LFqOttOJOtxy07j7kghALF8zLbcDiKJP
4NvSwXcd3vxINBMNx298oRF7n2GOfFInx7C4J/IogZohZmFRk46vpVkU1u262IZCLYEqoz1/Izjf
RDi49oWjNR41+YU3qBOQI9bEZ4+nuORnvU81hEvgImJ7aCwk4y+cEL0SKRDjHKyaRtu0UNiM8B1k
m4Z9qcBWsAhxXJTPRTMPpT6z51SQ+bl/64Cy1Xm/3vE642iw0h04LfKYCCpg2Sg+34YPisdvW/ct
mJEHXg945mYEhhWdMcdEvn0lsgum0UxAZMWOr9EKoyagu+Qo7ECRNFC8kgVDHvmezfNmb6y87Cgt
eYW8AzNtXG2PRIwxHmffOKJGbLRzj1X361vnSzGlLMTzZOXnRwMBLbEL6eFjFEm2uzlVCAA2+CUS
Vm8QpCZw0VNqjDFz9ubMS389P7eGSpLBukHyAKElU8OgLxKlwR14u043SJrzTS1+osjn7KuOF4Gm
4jUjELr7Y8nxRGTc+gP8jstX5KXd6G/6wEPUaPJM0ZMbGxT9o5nkpEa+TtlVv0nAfhq+fxixm5i8
tIePDP5bDpwY5UgAIXDkous0E/tDAUVd8D8/w85NwKfGe8Dmmm2LpQW+7Vkzueuv6W1kAStR/xXE
fDprQE8y6TyfknrRdjrEhDWY17AvTUENDFFF1CwgyWDxy+DYZ3ANk2oy4sJw9jwrA1eOhU6biPcV
k8j9d3c039Bf5CLLTC4bmz/ciyHnkSYhEAL+nDP+QkGxyVZ8QdU7k2XitKfptTZYtKgb02tRERC2
M4b4RsVZDUnJVYDqCYBDrAd3rzqsbVwlTdPP9Nz5Mh6AUjiz2SL1wTHNRnSiUPeP0UfixSVjtUH3
sppC9KAelJb2gf8YYIlv7pQNG4yYQolb3Z3RhQVLDLXtpYIgO5ksP3QrmN/rpDaDFh5HV0k86oOb
i1N+NFe5eZ82UA4j02DD02Smu37fmfXh520uPT3ok1GaE1DjF43nIxvnhX2rJXd2SgnSKR1lIB4s
WwFg28f35MZi6yWNZYvjR6psLS80Z7syn4QWKM37mIXwv2IRKmC4WXaWVETRXhtkvmfkIzl9JDvj
agzAq6e3t2x/G6QKQU6S/vMqBDpgQq0TnHhXL1kxX+MnsFSuuUyzvhvoKRW6k+zJguVLZjRyFh57
X9yMOuD3Fcgb3ER7J1qPcPtCqT57iSYsT6r4J9ijwgFUaY4SVvsXMYRZA0TzsrtaKgx5mBYXa5bo
v/nYqqX54PCgPXV6YG5u5keiv75foSbnbF4hLQ3OV9PWhe5DXZthn5E+Usd7uLPhAZHKazFwYrCK
5abC3c6HQoBmn2iMMOsaI6VpnK6Y8zOGslst8UvvxJnaP5f5AeZtyrtWJcaN1sZlyqWq6Rei6ODE
yivjtnH+KLV7uk8SwkIciGX/6DTZiTY0rQTWlKCMQ+xneVbcuAqSthUBc1K+83nLOOwNl7ku3t/Y
TwAC3C1drpWJNEj9iEqpY1jxdNKeHTmc2Gfs2wJE8fdp7Ff7kJNYBTSHWyOStponuWKBuAJ3MDGY
dK8zVWHscfWATvkYqu5AXd2KSq6ispp4K2kQI8GW2u2owzAZsts1V4XBR1BgYDeNFBk7K+GIZ+Xe
iN0Yf3JrsRfinN2+EGzjJPz1HqPfH6UBx6B/RjaMaZeD8M13EpfD7srBGZci172/seK/3nIV/HwU
eKknWpd8EBZ3+thfHHEWy/sjLYucYKmLuMwSjIjcdkIyTIe28aiODD65mJ+FIQbE72gLHMgdVBPp
FvqVZ0Oicqg0RADBBnH5AV8SkD9/NjY98clceESrAOu5jw/orMh97inHZ1I9ZnIQwyZF8qfma4aK
LgGlCnOEvAuyiJmPvJ15Sdd3y5DP5QgS0WtiU0LMyYW9VrCW3jqMqa0pKp1e4Zh+tig1nUnvAkQ5
uy6mSUuWDyzmGgLpYk3zxCoYNkaW6oqxb3aW7iffeZXFeGJ6KUg2H7PvsbgVqPxSLiZVq5IAO2OI
n39JWHXliK8YtCw5WSoDFYQOQnjsdPcXZ7+1SpUmQvhXl5lUN3qMJtB3StBdj4HrxwxPy/NnVlVh
17o86+PO3ToR1hXuRrgtpriLAqvLkEplzLgTicXvFJ8aLokKnZvwQzLYMhMKkHUZbMOhTGSY0Bt0
Uo09k3RAL//ngjLxXpeF8kL+eKZ+b7NhJt2w9wM+gx2uHkrDC94iRYzuHcmK1L8i3d03nFXcBjPy
iW+YrhAcrgszPiCix4jX7CXRjPOB/Z/r+dYDD0teC4cKnX9hMQkjRIqB3WMXoRg/HBgKzqcZSTcT
uyoHzCHAMWJXwxWSG9Ok6ycziPb1KlGYdxwn7/agfR2hPhs/BT8xADrHze04GxFO3SZTs59+fUkx
aSOmuJ7YekI8qGIUGMOWZ+n95RBEu5J65+YrfV6zg1ZIzGmpImuEiXX+LVv5cNPp+eGNlQVxeAja
S/5lNVDt5IsZJHTXlegicAtAmmRH4KZWmz4UIk5ZFV/RyFdVkD7xFBWNNerJHnivkzgvDebCwE/w
Q4kDiXNd0uaclZCZLm0XaPmRejE/jEKzxq1eQDG9KAJ89qx7aYt6ia6gbgomvtEVs5thWpMXevWD
fgVB4ptsd67CKKF14L4ckMmeXc2jf8wncVJDHV9/s2yKhrjJtlKGIQPgrSYTBnjOD12EJ1/GZ39y
mZ8n/5mos6NOLe6h5GYLO2QwkRYKRAjSgn4YWFF7MN3BT66xp5aaG1wtLo9s3Ro2Wbe6sXEb5Wyc
1TqiAv5byjv+eA7IwNSDpi00bz2kMp8INsc2jBA4ax7meJHeQm1eZUraaU1nmZQJTzcyNS4QsLJn
y9Q6PDFURMExEzDHk9UVAZbTCz4Wkg01I84hZqcqrOLhcyNRAdWq0Ygn5OMvDaQKzJbI/b8E+xT3
iL8/w/az2ZfPaDhWjBZZ4oSsG+pEZfXpyC2ruRQGopkxBrikyhaCT3omsRlcj9aR5hRtOS8YK2qq
Ijon9yyqGNLaUz50n3Ed1v4YE1+7VKHrDO4+cwr6BZ/OBIuDiS1rcb/6LuRNy+eaZjETP4gdnxDq
8lnru/O4GWfOCeFdyN1n+J+uj5vx7ukK55R5n36yAtBKSZDWITO86vqr/GB6a8WRA+CDyyvZGpTO
hfSWl9Dq3e2JfSAPbdy5lm5skcCBTnzCnbn3LN1fyAKTLykGFMoYrVj7oo4c5bm7VevWS9MJ6TCn
gJ2ByMJwwl9jbyAm0mN87pqcNPbuYvq7g0xeaY7iyjm3W/Q6I/cuYm4mkiNxBqfoQYK4ob0wIrod
hDqs2Dz8MvY0Jc6bfhlFgzTXbnXY6FxcVPkkRw9xcN/MSTHV8Cw3fjcJRSxzbAZADUvFVeouTWrW
MM0RzJdblHDPyBMPjpTZe8CVF3qgWxS9lVz6PuvTfRu9QzTmtoY9HfXNKVrMuwo/H8Z8X5magVVN
JGjAv4Lkl42jEFG2UkLq9xTNFY0UWKTyoRjTyKGyFwWJF52UH7ky9dAkWyL3EXUZZ/GYD8D4Q7W6
LHdLVMzOwfbuFD23vHi3RrOnoWD/jX5V+6od+LNsaMTVhWHKqdfvE8/3rs4o1zy+Q7DU/v1d+urf
tv2l8Y66n3/Q623aUNnukaCbS5nc69soxwv/g3pl5nph9cWEbTKepEcwlyN8GClNpVgoViB9TQKb
Ge9cNJZYxE88tdp8zLIHig5KsJEfDyFQkhIYPKpUZ3EnO5GsWU5JFh3EXtHkWRGo73ajAewaaD1H
UatQBARNM/S1JrIbkLf6dZk4hU0jihwX5s5Ryx7DNiWWUR6VT6ZpaJyxE95GwhomKw+v7hMnD7mv
PmUf9W02sweabjCf40TIWaI8qHSsRbt7islhI3JwQtKaxB3lF3cgYVGD/SPe3CR9fXEhGfxiHtVm
y1kKBak1nULKNZhenT2/NqqjmAn1kO90MftSEv/o0V9Erpr1fUI7oenalNgPNbm1EkCj0rkh11RD
tYsp3XQf2JzBJE4J4ttYTYFgw9NrjG/Jg+i5xxzv1jmg/fcpNV3fpJZBE6Vwdwjn7N6FJoDWG1gR
GdJZr01JTDsKiMV0DZOqhkfvh0VQDbz/Kc4aUtGMPTFDzsy205vrUlZqONKpVcrBEA+MUuV2p3XE
Fz2yzOvLKUSS78+PftVM6wLOhNuQxmNhVpbdx0vXKNnjPUWRwuyvG3T12Mc0nC1u/X1nKFfEfxmT
fV89aI4GfKNVaImREyGJcBaqxr+e3H320VhxXKem38D8zMo92X+TRWAcIHVxMkyCRWyvjehfX7gY
0riv7pEO2SRc6iQH61SJGS6vrMpraypBDuXiHlr1IVIbMFaVh4RhmKBXxSq8fPM/BGaujVKQRFGv
hWn6CNAh8XrwLTNaFQTFhREkwMImU8FFBd5JX2H3h2xTRzVsdnk8kxG9jZtDm/H1Rr2kZyOxnQ64
vqV9hQ8m7u08hOSrRrCf2VMApc201ptTbnxc3eXG2hAcqq2FunFQc5c04MeNFlkvHjtQQZJaVXnQ
VfnWTdXgozPcx4unQF7/WPA8yDYKa+0A8I0ByItudCtLT63mcGJOc37FIKEdnvpiCM6x8ZmswcvQ
BrbHTgDgS2dnPySy5WdzV1D0qow+4IUtvv/1Q8bbIK2LhJCZsfS3o8ZLqrcOmwGeyxuOor3vwjlj
5TDAQd4uNB18+Sd3zNH2CCDDBwqf4f/GSRmz8Kd+FXKovpCT7CseG841F9x/l83WQGh/IZIp8eya
8HARotIv3Wi3EzkHLIbHpm7aarKyM8oa9w8e8Lg6Ps0pjDDYUGSkTPeK0t8z59MBkO/uJuypTDu/
x16pToVeITceDaK/zY3wWbjMMj/qVVsW+7uA8ncDfVB7RXNe0msuzY6HQ7PKY3M5Eql7UZ8gzYZu
BG0RPBzhmiiFoey1m/KKpfWzKxUZisRkh2yOR+CVIQzjYbydMRXc8XJmz8qDU6bME51pLxuBz7iA
vtrucBjZZwIMb03khQvXsBO4nTHP2t2M1uNXxyi5aiLvx8/j/9LWQSVXtH4a/YKCtQ44jgWK7Ozo
jihb868MBnSq4B+fohJtP8ZHJvfNx5k89i0WYHUawukGbodh7542+YuRsO5FfslYijn86g6J2HzQ
/gf5KjY1rWxcZs87szspKS5vKCrnYBdXdCUxK+TQtNN5eZW85K+v2O9UfenaE2vzHobu3avvufEo
xAluDmTMOBcW1bmruwcnj0CLWQdKtAldlY3SQNquMPAFRcvYk+Mbz7Ofhe4m9/S6K2tEUBrdFzOl
yf0gUwAHyo0qXcZJr65wJVTAtsM0aJ1wKRuBeF56aP3Yx9TBu5czaloB0H+LvTtY6N7p4bK+6kHe
QWP7gZ2ERRKhwKm6l7Jdqh7bKpGiMTNzMwspqM7BqFqF549OeN1Gskyld/pON7mrEm3SwQj0I3ZY
wVXVa4Zo+AfKp4cGFKpFCvQcSPYKdyjsalXYfKf3fg9KmOc4/XOIw4LVdN3wcf4uUcfmR/GR/eFa
4qyrb4/RciGotkuxP5owzBBZyKyOT6app/ecp3+KhToNfzfvj1e/MKtI0Wm6K8A5nqEZHP0RGJAj
RqREf3yoDMXoBnEkyE0anPro1lo6qGIYuOuIPcP2h7lwJocdv9NPsx64AqiL1JaE+lgh3mlmVFuh
76DT5CWGvkPU1HweoqcZDIAJMJN6ZjMAmu1K5DvYzL/pEgw+wkuj8yxijb0a7KXXO5VjfBcyxYyV
NOL3BaRuhzz2/pqp029g7W16iDT6GRX6QHV8FX+g4FL7NnLVJ59kQKiKLj85e/C9Wz4RL37+nYbf
kRDj3/O7TtDfJplmRyxUQk5D58IziC1i3bTOOVM/fmci7ZEflgVbget7bBfBLEzchhNQbIf4B0uD
HsbmcVr9eB598TRyvp3xqD23ADK/LtsvLzOWzyVXQUbrPijrpBHVygV7rGXt2zDO/iM+LbIWK+6J
mGt+hx0J0h5GVPb4li4NIfo+mo/aSZp6wyo3PHIdSR9U/1EybSrGGDYAUrVO1lQt+WtaOZhAEZGS
bwZ8lrhNINq06PpVc3sE4EvRKPNMQGlQ+79DIkA0MUPXcFrRNydH2bkLVeDXqGE4+JlI0Fz5oL7a
4d2ovM6xhV9/zDog84l3Ql6OHV40rxEcKu15cRPRXtqj/hD+F1xJuyzbwe3/RUsES3rYM7UIvTQO
OJYKD22QgWuz5EMSP88Dg2TeAjS3yTc+iXnhnL5AzgaimDxwljAcA+Cbzi8uwnXy2IfylIq4Mvwv
aSSLialuUHmu78sl+nL7LJf/deYV8f3/fVpFtfx8pxwVLpoCCJmJWQQ0XDeKU333bvTtAaw2tQBc
wc0hJJGwiBikU0WY6W+K251A78Lm3U+IR7uvEECp2MiR71pK1mFviL2RMynGUCSSiv8Qo1S4muR9
O3cf665wuW1g5+KTzycs5A19fi07q0M3ET+KgMqI9809TBk3HxDrXHizobh+r+QHOUDkxHRYAyEg
eq1lfOeNp//TNZX5b92Zh3Nj4O41tRNGlRTS2i1UGfoYoorajhVVom3uEdYZAl313Tsl8DWBQ8lV
j54lQIKjERSHodboHNDSqxMd1vh/sIpiSBr6Bw1uoR+dtriWELoJP2JvcsAOA7/1ENHZdswr0/Sk
i7hCI8JKcdJ+bL7YjzE7WIwySRtsPP6qDrDr0QyGHvL3VgcOWD3VgyvVzstvJIijxsCVjmid5B4k
7dwrEsZiAepqkIatStbFyawvD3jS9An3GGhOTN29Y0EaP05jp85+96+SNxABbXmhRORFcR0fCrNW
XHCSbqPVuxGFO4k/xc6QOI2d85pozZ9DcH9vgGlog/7/PTefnKWAYhiUILsKhQKoKeacW1A2VnNW
E25Xc4Cgc7bjysdcAvxh9oiHw/ZG80B0E8AgbfGkxB3d9agykerfoeuBSgOGyZkZnFYCVOgdeAjG
2uTNyVwnZTtsoqwfk+uA80eOVH6yv19DZje5Wt8SJBbjjTepSSs1xVT9EZTek9PHoucEioYbPOqL
e39pBsbi1HznNEKmF8vZcoNsI732DOGyxWeuBya3BwmM1ot3RDhGdv5THR9SpmJNywczgcf26MJy
5q6MUc3DxG4z6ZotshMRmh9iaJDtVyKvSD+BgAxY86HRqpCR1k325yMqlDhuoNZRYrcGk5wQYCud
h6gGHRjSZXd0MoMnlcpXJZ1w1QV3L5WvDTVHPZol1YBFH698PcHwkAsasn1Po84i+jOpZiMaiNLi
DO6MQFMsmJTSsjMbULcXJWAmn2slh/5CjbdnJIxqEP0wPCPt/kULK6jsegC7ZpUrDc0nvtbJzrLz
kZp7TgUSoI3DFimViPuPJtX0iLlRoikolckeQgm9JgYQ3EEuIRy7rhcz6alKPfOd/fN1shx9HxR9
DoS4uQ2U4qXICs5pSeUmwjQxUvK/vdMka76Oc/TvaYNHZx7T7oaaXQ3q2SdTralNDtnzp90A3IB5
dz9BQke8V75b7jy6rXWpkC3UzKN1dqRTI8DLft2MLDZCTiWwAB9rCv4FfP1cXxaPzB3b4BGLTR9+
+B1O8Qst9Qn0FELhVs87iZcQ2nVFIj1zlTRRWFr/58SgecJ1JnPBhKuCVpXkbdeteOkUj7s/1gU5
fX1QNE1aWQYkKLH//dZvqBG8NwCyQIejPf6kWVvNqR0dM3ZJ3MUXg9Gsvm6KrpFLKrtn/scO56iq
5/Kdu6hEdfgbSSQUfy0iOJFj40sOn5Gs06DDT1WLqIP9rWM1oFqxjYV5DtnTrOEDAx9NhONjH5cl
jibNRttp4CfL2N1BY9PfGsgdYzDklEupPl9zN3k89ie+4x6u2v61Dy2LT0j/mP+I/kTK6hRobLdS
7oeKOUW2st0xEOXwpK0L4OE0H95n9fd49iZBXTQ6AL/CI2fQRHyGZVxfuZsDEHqCKRv2tuaSEp35
dz1OgFmuISUygZiZiupiqatQsAfTHfWgcoVBiq58zoga8u19mRYuXXAuWVKovhyvERADQxSuw2xk
XA7gOkm4JKIftzRFpsGduSby4bIIQKAmIg/qTLhqi/xAqlnVEGfOBHQFnSmXfJeg0wI91MHXlZGP
VQ8iZbn5G8KrIXjzXBJ7HDewEO5V9mcq2UZhTxk6ULrToGd/dX35PAVSax3hJGpa/edKyu/MR5Ic
HHin6P+RboP5aUSlaoS+2OfDagUvQGfDRszWoV4N8PxjK44qqRfjx7ZZTuveoK3cix4xMBh/zDVl
D24MKoSIyQmYkvR8XzgUkzvNHu2JNafaeiHGAh4ufsG1Hq4+LtMTiB1RMKTUfMpbwp+BUavZUHOh
vfo3erkII4SHhVLEMwlmVE0jK2Er2WffjG+Vx6WNtxGjoKISRQtDQkGkHygH9QEzv1c7DL4ufw3j
5FNvy3EXtnVvrfurcn3VLIZWHrB5/d8G0crIrUBOi8nVodX7vIV3Lt9OyueFgq3R3s2d9m6eIEv2
8eStUI2LWIyBglqFaMQfj4dDCliekW2TZDeg4SDhGnad562eOOoUzeX682/+ovsuQGT3KxbPVvhm
8UquO60OzI1dmW3vYFqj+YwX+x2GtbsamB7bD/oKRGtQCvYH05PRHlskcOkZ9eOAFmoQohrQoKeu
hqWa73xx5hPwGC3NiTrKWuyTOvQA0QmfVXNqTWhw6iK5e6bWsTX6I4O/3cL53UiQw9+lO/uiLpfy
Tc4P/Bt524PiTYmc6/rjeZO5GRAL2lw4uAyJNDKhzqde9z++Hr7ywvgFtuEFRU7sdUgBqjvUPlNS
nmvZblHKYF1vlJee70+G6zB7u1zK7CyqKyQWVNv78AwjrDPchBupeGkvwMmwhenq0OX8GOD+McHR
JJl0bNVmuty0Bk+cvmy0jrsrgJT1DDJjOeLzi4YGIFXCd3wgRcj/HYsHP40Gv4qncNiAvHo31iqA
XqrD07RdkVzoznsDXL6erTdoxeelZJmAxVv0bnSeJXhhnosYV3HF1LypxpUoTxplofIPfuQRtLZK
K59KuaQK32Kz46Y84e9AxTNvTcsZMsbNptNsHLEgv6UcREGsoQIZZMe9fnmMrl7Rt5YylxWzfnYW
dha23aPikCsQKOYyEVAZfEhL24s9ICabraj5HPnpbCYx0G+3x3LqchO3d17qLCUKG3Yh0J5HcZnA
AwcTY82h4WEw9TCl/BcZfm502zHBl1hVVnWn9WsGZad+Nu2aKxo0O1Cead4Du4ca95kAzqJdHW0G
IocsQOeyMug+e6TamQu8nBbkmL0TiWWBZs8bMa2pk9/6OWyr+HOqIL7nP2I6wLklOvbz+LjhdGpK
SebmVfkjkJ6+QgGKJA/hKH42ArEzHFxodfSaXwjpE5a244EiB80kDsVQi8vJF4FKaApOEFpYL0WE
jQupwccV1IltkSQoGYm9NV4Tg0rpgPd+V/pzg+F9rcRIfMZogJfv/L5lqapgV+TzwE6b1x+BTxTh
A9m+Vg05xU2yYbiyUvGG2emvvzf127j7ux2wMiWA5QlmaIQOp4i9oxZ8k2P4HQNDtxhK2qSnO89Y
0HRl9C/rqoLa+MGD2OzT0Y3RMNc9HFfAX61DLtGvgjxFFkCReneRsNCqoXnGvjhNdZlrC3LCGIum
DmuABezE6vrfVus/TDi+vOkaLsJU9dLHAABbpWIUS1Coy1iAW93VRe7EY/sFbDvZMJ7t9DeQdU4b
NUKMNagYJ9TQ5fR8FUXvumI8VVon+5SuN4M0wqEDqbUbtYyOddMHwBAmMVoib0ByF89wATlszUhx
6rNzaEM4+tSscr0Bfs2Y3fN40EO77RI8DLkpK837HVO9ByqQyTTDAlFKgyjoOjaHtyfuY0QAdoLn
Pnb+PFhqbzXvuGlJ/SjiTIpne/9IDqJKlrdtGH0yx4CotMSKZRecTKyHmtRrKPcXy1cGaGQfhGJv
g4plzfdLJl5ZG0lkdpaB+8rdUeE4nZBIPamzkRcVbHM1SvIb37ErZU2nYNtDt8s0QvNLn8LSdH7b
C5SdD6vhVO1tgzHHqs3d3LvzYTjcVd6mepLdU3aDYAs0qsroGpBQvZ9zwE/gi4G+7l/nt24uvfAk
KXKuef6U2xOyqoTPhWONgBNn5qPtm2bdnB02Ozcuoncl0Gp+58FUHlX40lPw1nfd/KEwOeLIKp3B
mrSxtBYnhOYYmtjeZxp8ScgOq/F188nAazqlvtmMSpB/W3MdzQHvQ7MoxZeP8LsipieHWa8aS/yZ
3lk6+NmkZreL24UhQdVMRZGl5cCRiwBA3BSZudJTSlupA9TmpkGodLjX2RfbaBMSj+7SVH2pko1N
7xjVMDfJkqEf6JJvBp9qOs3cjXS73QhC4c9MDB5LC96YwkROAWc3K1AdEFjZ93AjkniROgPzNZD9
QKZU/iIfg5oINWmckZkW1PduxoVmdBH+TnxfWPHInhGvXWKNOg45mkuM5yvsbtHN5yLhGnLzGk6V
6jbhrZnctAhWMkCw5SffuNA6GhwW8QaxXRBUd24YFIEX9o0JvTXLOJi5RYg9cDwXITpILtk+3qJc
5b88T24Nu3a9fYaS0VCvwxGPkAxiMY7z1GTWrvNwNb/07wgYVwC8gVpQy4IELpXJNt4iQ1TGwG8S
N8MHVhga4tFqYQ/yq3JShRjJB6GsxNADB6j7g0Vdwa2CCMYBE0IHOYvnTom3fgWQlMtV+dHVTEo7
fqcyZf1jflEFI0p9gLU5qMEg/DL6KIwcNGku2FERcbppHjcED6rOAkQlyE6twJ+rLgFEIW/VzqzK
78dYpQIXFIT0WM6yt2mwCIWY8T4DqDv1sl1nbVV6qwakJaQWHL1akmA9FB/T1Zv5NDRRWXDKQsCd
fmqOlQOFqeXEoeUaBw72cb9RU34Qc8WNHIYhq0obqk+xXwsMCO6HcDZIIiAKuUVKwTcTEsUGCwhu
EktmtJcykVQxg1xaYiCGsZgsrwklyjvbhd4NF+XWeov3+qu4fpkORRmaexoQICrpMSEfOSxSsl+U
fKrJRuPSYXImvfLWdirGkK3ZgdRCQWa0UnRe5DlTwEH1CzrGKp6/FoT1RvZOv3Kq7nAxyfUCEqIb
nDyMScNQECC+r9V++cG7mQOh61H3Cp90axZOEDF98EW2tLdkXVhht+Scf/mYQrrTRJOuJWynmCzn
ofYmK+UgsQ5h0UXHiwXwdfnxoMAIE/0JXfXxaUmKveiFdXsnDrXWmkSkblEsZgYkKJgdKTQRLb52
IApY4BavW/oG2aLMLnUHyYz0b7eXbscZbhhWChkWb+G36KB17NBgsSVsXQibmRam/wYP9URxBrSG
OMfCjUXPOcEt5oNQ9Ge8X6XVITLg9DvnrusOC9NIH9FkqLUAGlAS9+ebwu+F4L3bKcrrLKLo4MDt
/2f48cnKntK+AoGVDp3Vhkc/dpBPH2nYQmpRREre71DHJJIChfEYdq0FrLLPAnByh7SXmPLhDJFt
391LdA1c8BStPc4RW2DDZ3HKRJ8eam03cnyDeDui2glMV1pxMoNBk1YyO+P3QG53bRVqebJB6rkc
88cgxuOY4KG8ow3KvSeFhlXngbN6GfNScdMMH+kQJC81EAEE4GIj+rfQjiobeCPkwnLnxX17C0Js
tmOR5cTACySWSOS6r6mgT8nD1yfAsN0UKsx27GDcoZD6QmAeUbPRhP9GzdtSNVU4Uz82QYGBCVAt
SlwCM0V4GjVJ9xoVjunpDuwojJ/8Ef5S9j9ZmaxR5qcz26sz8Wk3+uN9tX5sifSDTIP4a+HSAElf
OLyBPLeclv99KK5J0QtXkQh3tVfPlJ9RBa4CwIdUw8Jf2SoMnPDFO0gN4cNTyNljsrz0g8dJN5q3
clikdMadSw4SICl5faFok817LZ320ifoQvnpNd5qVeuFQx4Ks4KPYB+bvdByP/04ukd0QblDXCBW
6DjhRxrrTk0CgyhvmtIJ5Y2hsaLqjkPsSjhVKQGuR4hQXdRT7vtSAr3hh8PjvvGItZBJICd4UXmg
+dYr8tjvrAqUH6Ay92S1/FAA45AYyauo4C7D/Np7WVnzVlWnarpbaBF01mZdkWmtlbEkO2IjO0ag
ablLoPLXr9gAqnxis3OmQMZbKhix0bgu7Go4AMQgZueHhQ12WzPyvNfYj/WfRkuj64XMK1v1Xp1f
XF9TWhGJ9VwGumqC1FDquoeiLc6eLn0Gc+gFZ3H5WCxbkniolcgd8bMA4P8JAIpsjRF/RuVtmC0E
uFvDJ16U0jnETiJBdQ9c6KNUOgEUZLN9DEZSxyAUBMGb6es2Et5p0m/nTmefRuuxkRoWBdGv+e7Z
g1OxKqJioAkBDD58aDIhjeT+m/kcg5zoetV5p7+eDSSmr8Fg8+lMZjBh3YGobLjQAKdZL+Hf3a1J
BKyNFE1l2+sLEZGATJfsWQLKwfFfE4MUzmP2Pox8sWf7LOs9YrbZXxBPEg8lEprtpbGEOCf248YW
PuXkcUsVWKMGLBMyLUwAy3F2ztFrAEaDQt+Hb1Q5SsM2hqVbNBGU59Ke6H29tN1y3t84+i5gcx3T
gXyrfXM3p9nqhz0926lBgF9BE3STBDDjJidlozRxnmJjuSp5rF3kxK/JzoFtzX7aud/RkZKczrFT
wUYe4z5G5IybsNcwwbdBEvB+xmvk0X0trsDtHcCxf0CxjqHE5MkLVfO5k/KKEvS8UEt679U9AT55
HUJFDBYuWy/jx7hZMeZDgej5bdReA5qFpRo7fKeYEifl2Rt2/+ejBqbErnW4vNZXgsilwtRQxq8R
501yhAZwkFuX+Yj7jNXURFPyz+B/Yexn4esZ2HQG0BuXw13ZbXo62wiBNb6kX+occ7kKIOA4JYyH
z5qzM0Up7eMCjixqCc0HRrz2DEJODlZ2WVysgMwS6EpTkCvRBx3fHw1uMYTyGwDJ4ITZuGVgh/F7
dgGTQlWZKsg+XO7GYuTrWmR7M7qkVmWMUIm8YM37Dc5Ve8ax6/ONqL/9ndsNUvIXfiD4fFDghTwI
+BGaiMiqZ/mOsskXhuvrORVGEYK2sWTwSfLecQK6Zc9RvJvVtxifRuaCZxPKus9/prHlbMEN5VYX
UQ2JbctGvSaGICTIkqS53w43NtWJ0wj2cQDsAW9PnC4lMK5U0X4yxXMG4n2lW2Qx1U8oNmkanmzJ
e2ZEpGCwPKGUAHmo5BC/Mf6cmMnYqd/CFp/TGHwFt3axyhC3ZJxSmFFkWKaLUVmU/0x7mUEWPaZ/
OTnuozkJS5VM1O+Pc0NHmPtkAqo4PQkAew4srY3kyVCfnSiZCZ37h2OBqAumnD0xOqeIU6FPE9tL
9K+jnu46oL+WrfLqoWmzyRH3x456qIQt/kUM2Ph3Q/BCQCPxqLUQ1LuIleQ7F9zNOXdR4JfJ89cb
OT+QSDwJ3/OKGt41NuAvKL0JDJTELN4NnlMU8i2m6uJ3ruDJcZz9tuxPyzlWdVe9PvU9sZOTy7Xk
iYBiqsRYQDcxSB+T/BtIZ/YuNZtLeZESB1jsb1X2Oz+zhbGIMz2lIKu9TxX0WOQHCGnwlWXR2zBj
LdbISOvrCKr9N7yYYCJtGXd+g+stC30iCk4Je+ip1almA7xIQltF0sGnfp0mbdXmBWP+guNyO6II
yLayrt1840Np4g3NXlImnJWiCqbUURFqqcaBjJEO4nhPDlDkBvEItSY9NO0wWHUQPB+t3e9abGYI
etPQiP+ansr3TICI6yakk9da5tTRWRiIIe9IkgW0qlYDSPCwQ6gakjRdYWe4GBKVVykVpdeprThB
D4ZZ70wwxSaw24ysOcHeTrhrCYEy/jGUQAgVuBO/JeW0k72+zb7oad2YLHAbeiSyP1nclb4Fxq+e
WkPayBVdVDKsfjTa03nttCTdDXc9O3RoYec9z9XtwBq0ROnpDXhmzT1dUtQDWefO2VWAVCVTB5JJ
w21RnFmXVjEzJbHNOt44QRzEesCVMN7jAFQz/YCzB/RAOfpv8c1A9LcGavPc/87fwE5jqeS+ltQi
beELTK2rSvt1sf36ih8Z3iD/h8frCMl+mA9tytMimPGq+2wzmCdWIoVH02v4oGRfkjDTkY/CjM8q
b8pBr3PkUXf53GUPh9RrtcElKW1wtFQBx9Q7xU3AwI6CsekvyprBdUp2P07UQ6sU4NjXvyvGgiyZ
v/4Vw61kToIAsFrj2NcRQSbl3DGJ9lUK3bvexl4ey1LIDGQ26NaYs+4GKUo2ZL9r6CJh4imnxqqy
PbTlRrPMPeiuQxrK29tecQIfxmkRySJQb/CWFgtAoQ1wiu99xf0hsWGwQO+V29V9MfSwlQPQ/ADX
ugYCHBqZ+zZQWxWLhS4iLxLEGfFSLQp/tHEzrZ9wk5t/9AocF/GVxE0k0gngOVK70laGcLgbtvFa
zzSz3BGBGAp66+FrwKji+iSIeOpwMJs9oHdPwQe+ueABA7hJEzjRUpeVoHIzepe0AvWPeEndtHMr
WpwSEbNDQe6xve3Mv/4bA0gnRBdyoqPQcUkbDtXLArstLBoeIGwxeU18w6ghmQ7ptADMdDih51yI
UCh66ebyjDkxIjlcN0V0mjItu3keSYAaPkaZHi1w6QfP47rn0KdWa+qvhKW1TATnabLEhWViBYb+
uOZopl0S5k9KL30/HZVRvE1Z8MBHB+sw+z9jnHL57lr5IMXOn9CLYxmpsxvXkp3ZuUGDXVRaWnXd
EhqS0hV1SHKgbGCJDtsP2n1Fovl53yoRWuojzCPXlPPvcB+wBNpT49iMurgP0sOJf+2WoqlMeyCs
rGY8lEB4kjl+p/ldbCgM+4e3cpqeKRsn66utGS5Sk8ABGXPQJu2YkxA8kd/qP7Xauiv/8mZWqn9H
iygID5MzcXqjnruS36TNCp66h6BxddZFtY7TPz6WtmwkVcud3qqY3QRla0/DV7AyKWOD8xMB5wPr
CBmqfg7JG1SAtgGOJFkOWEFvhib0fXIwqFXF+RaMAVyhUespuDMFxG0BnKf4X0CSYPYcwfhij6QE
CRHysUFPUhoorjmi/ATzI1MqLwUDuDy/HYUnjwQs/A3J2f5TfIgMdNSBf99olUFFDzMEb8C3Uypm
S7V+kKZxsuOXvALcIrlImhpZHuQTZv0+BbV/pQw/5NtL4AH83vqXrhtSV4w1wjwx0sEDJfqkyTTC
MJQhJfceh4UsqiOSKZ0jiSE+GJ/HUdoh+f0dv/YNyS8Wklwj6C7/vo6PNQj/1U0tI6PKM+44+tKT
so0td4cgqt/P3e7vbTvAhhFUOLubyf/oayx4+S5SZse3f00tcWQ9H9jxVxdTG3YGbtnHMlKPsvBI
EB8uKzAybHNRGT/qka80YM2VZxIjJTSHEHvlzBHK4YpHdro+Ft9EYFpjW3fv+jjvQzYA6Ct9+3ds
kp2zE+dw7XJenInja7+RM/EQ7J7LRwqteoYJfAu6crO7fmEiGQ9amCLHfC8AhemZlXqks58FSZoR
e8hvFGl5wxnsp1YQzHY6Fov893Q3UYi9bAWhZRvkVU6fZmutoz8gpVJJTRbM7+4UkEnHNSFcHwax
6D9qCITmuXA06xlj13TD0Xi3GoMNtZYo2+LRaKx7r4eQihPejTyhFW+rouxaQ9v1B0Lofa+PsP31
svSdTSXEc9IFLu/bUR/9IxAlL8ZLlM01C1CijOtlS5W5aFfdldxLqtgtz2yqIcVli8b/XNcxs0+W
Ih4YJfoLIv+w9YHzBhAOC9+DI4lYRQwmY0B0eqnEwv32daQ2/rM3MkP+1QYpWD4x9DkcRPGcB/Kz
ZPqTdQsrHVQz47ogeqI2YF2Wrc9bMX6uq0NnA8I0VnC52u26mwUxKYueWnQcqVSoZ21SVs2/9VA2
7h+lfr0YipUoPRgyGGWTppRdqsAdhEVsTZr19TdxNq3LT4v2y0aQGAb/ncBEnqrQt6f8Zuvc34i/
iCb91RLjk2+Go/U/2DR62jU0D4DegyTblAL+21xL8+LLNBfbUburKAeSJ6Yzl03aj0XmQXvqOt7k
pxwtH/r8egeZe0WIeP6qDEkPLKkBGYwS5113TDtrYFMSCQ8GOz01RQQFJnWWOuMEC5a1uC5eYYy0
KB3nDPk51sg3H/VOy7ih19OIydZDZ6J4/RLtsQyz5Xly8I0dNC2wuFo7lHFt9h8Ex3V82qOXAn8m
R+WeYR4f6drQ7WWfxQxzOVRPZe4QrLwlFEpHLJAUyLi0/jYpuHvJSfg3jCMNtHKnTOuxdKbqoYua
zlIUg72up9z+8TWOJLKv1A2a7B9zydSumo97sLjEGK7/uuA7pr1FR47Rc8UyroAHszzGjqe4usyv
CPZr6yjryccqReesO3/imDVJdLzOu2Isgv1/HXE+pWRKlimqX6N+R8Mci7IN04kyKjoLqURO4rBY
GL2E1DqJjlcdY8hMTM7/C0GVkQ7+gsQWxPDoF+3Z4pv46jDztESk4aiqtm2SmepaDiG9+4e2BeEY
eeBGf/4LJkDbDvWb6B4WEW85qRTBgbZqZexmYghTjv9r3oVwK9h3zp/gYM1SJQ8noB+6H+GJqiZ4
ht1ytgHmZ4+SsZ49yVrMrURB07itJll76DmgNXTPzQ5/4DP33FHKmIInkVjlG5r8bnn6IDH22yvF
8/4MSIUAukTZbyey1NVgkwv8+BgNCQtq3ox06r6Sr9Qw3nMV+vC3/XYd/qlJa7LFsQ+XxH31pV4A
5xYIMPM/bSfhzSGKD0sfLnITOunIpabP6D5kAZO5dR6CRfRntr1s56y0SD18+qF54dfr7XisOHPc
7CBp0/s8f2/eTLFi2JgyRogaSByZVC6Yo8c/hGTSSivsjEVrEwcsq7nO2hDx9UgJ3azQIozWkkOR
inuQ01UP8k0PiCf/qNYANm/MkS+QqwK9SsChiTIqn4Hh5FFO1y0d0GTYyd+aRipe7VyN1V7M0Gn7
ygYzAMNXuycRO0y/SF2gFNuzX7ZecrmdzmUYki8JYwUKo3ISN+TB9Hug0apo75ZK6MZ/wmDDlGJe
Fc2rwHzm/l2l+Yb8azLorHwa8tmCOIN7YsGBBq0c00b5LdkmWClXmaXCFLtWb9AyGSsc+JKvfnEi
FNvcv5leC/6imH2o5kjPNuwKdnaeLtULuwFXQrEDCS+jqTMIu8hlSJWiDhi9msR6LmXsTBc7H2H3
BhYqGUk1OJcBEh5tv+CRssViUz6AFamaXcDJ8RtnqnzmJSnEKKVgNldpoMSUJ1qMbIflqkuD7ZlM
ny/FqaM2RxaRaAVsryjSl+vYnP8alGN4FCSxXIeJ9zYfL1UB5YYMWsuwZAKpC6JWZOLBmduNvkeO
E8s4qjFVeYXWiN4dwOTsU5waxfxglg02enZ7QBywgfHFt8c8f+zxKnv8v0E5ikska2C/OPOUb6se
cLzogCMFhGCQ+XDAEJw6VEDT/lhpbaxkXR8Q6kF0gk26wKTXbisYng2vSdssLNMPVUYjrvonBbsA
2V6NBRxNrzO2P0JC7TiJ73Cx0ka4pdV06wlgy4cgeWAj848V9aHuMC5UD8u5sBjufFEHjB6ddqei
uYvmChsuJTq+B++hobAxyTHF9j0xSCo3foS3EbeiIKqDCgIriEen8lchId0j4IeKQYH/aOW6O9/z
re1y75f7CbHAmhYBC1ohJL1i24erd2lb6MJqixOgzPQoncqjs3jGPYEbp1iF7mMmZ727CooSuOff
tgZAZvX5Pdd4y/0G6vu7I2w/b7CmlqO6MVU2ATJS9L6QrrruFTGlbbDtlzIbgzwOK9G3kUHfEW3q
GkfvizfHNftmHHUJIheWUXyDSoJBndade3GEa4RTafyU5GnxlMS5Dea0UY6C+IQksISi7VrQZoX4
LlXgoz7PJNChmHVqBCeU2YXTawFsfxyyJMpiZGuUTGgCbo5AoJeonKi8kApMNwdVTbr0IDMVdXqA
kWwJ3iS7HxUjuWQmj0dz2ghjAlhWkWdkVRMeNLFi2AsiBvbsstfgoNpLxP/tog9glGQgJ1I59kmM
kTdmsk+ZWOyXWvrP2qwcXh4/d+C1jpwUjC2pZj5dsDYRVqBlHhiMboz5w1uQNqxme9L6sM2+RjFt
mVwbQ6cKob9KdslgeF3yK0dwQ10jw7SkiN1aoWVzB4vibS/ACG75x3ed31m4kBDI4gu0AP9wUHkA
nUtv9+j4ao8HGjGWuQtrBA0LfteAj4+bA7mEj22ZxR5Z1xHVr19fHEpuaCHs6IbhtOuMr/NFG1JE
1fwLwcH4dnrkg6TduWfuRyV9qJqo+w9o5PfZlrkh7o6FfS/hvMTwiTHE4ol3jz2+2a3LbTJh7D+R
yaPVHmN3/hgEVwzzHe/dT+yQj13iYjHchT6EsbEMdCR4BgRd7f7Wzr5DxpCOTUGGolqLQD5Vij27
c/cOYr5o4ffxeR8GVzbhjxCYiDlY2gFCjAeaXcSlNDThEVN9SgMHS0iQtmfkvISa8DHEM2UyjgDV
PdZelfvdqVFXddLOHLybsFTlmIu1MS8Vx6Psq1b4qAvIHsU0V+QFgglTbZcrYqpXKUbgTeM62lPg
FURq7BgymQMYUJ5FXPJtHd533tJGNVngQIsyafMlJxwjrMF51bDaU4N7ZHNR929tNNZL7PSjEvXu
Jy9vzr+OV+2CIyAAJLI22lqcNzqQ2fw+AsOFSXuT/A1n9Tm6dNO0Twt2JI0AMfV2rpvrG4wXjl/S
fF8dN3lUegC3IGXDTiJX2l51S+OXlla64ruQPyvaH3JYz1WJfkMIAY1P9PoNEOKZHas3Tz9WEvwv
D0adzKYFiBi0ObnuK1DZW9mZcPXjYf2MRKLQVLgKgjOAVFiJPUQaZdL4VJHZaFhYldj7JqsZJXV4
9cLqx2uakL651BvzDOBDIGj3WRrUjJZeIpNhDKPtxSKjJs2k499FKn7z+/wMdOTdElmgqv2Tqw8A
apBikkalTGwU2ykoB/oJ0N7cg4dO6X/56Ac1ckQru9k3tEKiKEh9syimGmuLxSpwCLfhixGELR/Y
XnkLtOp3i8u7nZezLz6Ntf3FV/zrje3gWKm3BMe+khFv60lZtVudzNJlX4H47VVOSmtBEjyHlnEg
8S4eiCYOr3hBZ0vr68HAPFtN9k7vRblDSaMns9VlHq1O5weYmCXW8AkSL2b5fuEpOlHfcdlBulSM
F/bnV2IJ9zmmTMAWq+4xiW0rnN2Rln/JyZ3Yu5qfiAURxNdvVbWIdELBu8+dSzCcfZq0Xht6qvaR
KY1IsIROlTaLoFOGSQtMgvU1m4maXtxgTRZ4AkPu5wljMfpdrShkhjtllJf+jOr4obHgHVRcTnhl
A7E5czdFRSH2tELtnnQyFsHE/ITVlmpCe+Ro3uoAc1VYzwsw7Vzv6WrVZl23DAHOHQssc45FkOJQ
jxXISSO4u1toQRtumtn1tTJv1cNNgky8GpLcSAFpI1RQh5Il8Y5J0ZIMGNeLlJvpyvi6qGIKu625
fTfyWuB97VOmmx8+v470arU6CF1B5nURwTx8bphZEhKBS3GIC7+dJBPY4bWlVOuHyj+Au6wMhj2e
80gKJhk0TpY0w1cbZxvFy/ZRVFHzgH1IvhFboVdiiuLg6UxxWvQMYxxsVmNG8ih+XJOz9annqbcC
UCY0unQxfJH4kLVq4RqINn6159UedmER9PMYaW/k2mAKNNHqHWt4MJ5TIq5LmWhLRsLUHOiq5UQi
G2BffqQ3GwChARQm5kDXcM1mkxc2buNTqpWxNdyOWH/RCXmcHgv8k0gE1XB059JhXOq1g1DS/9J4
te9ZkE4WU5Yo+8EpgqbVQCO48AkVShvs60AimG9jPq8ShPw4jP0WNa4CTOg2Wrnv2U6fEBtWLgp3
Tc8hV3PVUGE+yqzNOl5Ud7giv5DUS8SZNO9QSOY3mr44IeXbUEATIyVmofWuSHyCLmC84H4nXDPH
PN8fVvQNKiKaxlo7Txf5pdM+zHyHFPpZymDOvnsSI2ZWRPx7siVXl9oBHFiyiWWmIt6gKD8Ox2uR
pVEKZs0xThQs40kHXbDGXXcTgErxx3qDi2obL5fcXbbALhZMDcqD+OvRMpECgGKNeJlzNOUWiI5H
6qpBEJeM/yEdjSS7O/46oRQCgbqEE5r5LlQpnuH7METAVG732dDhrrSroo/aNqA4PjLmiRhkEVgD
b84pdo0MH3Xb7Rmbi5diEPERDWOaZ3Qr+diXjZbkpQwaKQwbpoawhLJNZ5IjEKFsGiFKqv0nmHv/
PCvAXnoJTXLrz+dooiUIbYNF7JeMhP628GsSl/+pSeAxVaIsCdQr+RgJSzUVe6jJ57vibEilNzPC
uIhjO1ReLdk2IsYXI0EfIJh2IsnIk9Wf+UDb30Fi6OShIm+LrbdnUH0bRjk3BgM13oK31dFr5EAF
eyv2MZAF/vXZmMTNELR5MDZs/OifPbaV1ULX6eOMgyq863/Ovr7QPziaNZ9oxJtnjjgUrrtL6eOr
vJq30/W4q5GM0X0aDFtihZDMeIo4VI1G9Tr39cDkYGEgdL+c8L6HG5QcDKqV1QJ3a0JR6frANuX6
t9OOMJ2WwPAORGDI23l7iAT99gjzGQG6+6z4VC/mvSUN+lNulZHRC8mbC/g8WyR8/PWhMLxzXGKy
UeUCd22oHrW8bIQJrRnXo23gREWcs08H2bVYKigvLSKhMjKx74VP5nU16T5LkgNvNk9wQ5HU54Ou
EAu6VopHCUcsz4ZM4QYHlE2V/pOmpZQ+pQezgDVRb9Wt7bd4OSfpfK6kpMXm/gNP9vE1Ts8VXCkM
QH58lRfArGiLAisB4maG5Z+d94hpgMADmB6HJBve+xuvMY6XrG7gqsvRS893jvUZfycKe4EXls+H
9VcOnnaEVY2sAHpNJfk4KDwtciij1wvXh1Oe4tH/d4Bs7r+v3CpRNRwtZZVDCkSfz25LW0buCuVH
yqbOXX6+1S4HzTXqSLvxnxN3Xlg4LskNwUqL+MNg2goaEkSXgNizzfm7lCdbCq1yYmqDJR6GFQ4B
jNZB2y/Y3jCAUmSw/OfVV7xaPa+1bbSYj1Xe/ev9W74iR21pBHVD3CXPdu8NtlJtjrfmZpd1YEWL
8kQxL+Pqk1Re5G5vy3mv6LqHKzIPXHNbBrxpm+80wlC7Ms+NIVE8B1jhrVmMnZksOjttUC3NtEJ+
zBQKrR4ndRDiVeCOeM8MAwxHfBQ4LoP8vj8AHmI23dlUnbhqVUnm+XOzZZhhvu6BYrC2bttcZVXU
wreWl0j5/XMt+ceo7BRjnHZONBl2XFvPsApBga+0JNR21nixtEt73AG7a7eTt4WRGCucQn0scAbU
q1ETA95BBMXfaPvQAe1UdD1PzQdvwDHcXo1oCZ0XLeYZ2VyBZsaARKrVswqbaOx/jDM/DwRLE6oS
xoNXFCbtWYx5w5klPjagmSkgvp9uRcG7FJnQdgv/WODkabuwKW3UNpENavfB7frCH7cwyJhQUS3z
iOtNp4rZ7pyOq9+7pubvUaKf8fI4S8a92zvSXArWFkx3ya57AlD6gGJ65GQIr34HSYb0lTj30JN5
YgA6PzNvORsdlmkvqnZ2l4O02jpbmfIPxfWoJ/xUwHDztFnYdrqTpOGVhIzlqHmQjCBGT3XmDYjj
tWgvfImzYFW4LIyizV0LLTV553O4g58UJkUykUGjSYSVbhFG0dAM57UXzHgN11RZowK27Jqn7ISq
HrSc3iyZasnl6CtVm+g2/YtEWjWQ/ngbPlc7unvRnE8QYssSJa4hbsQ8fmE/d4UVhh1ef16vu3cW
upVXsX57GSaCSZ2FgG2sfhKEVxHyVWtgkK3EnX6ZUufaE+LLKbRzGkrqTl4irMG8vzreHZ4vYG/4
Xy+OsaA0iZa1FdEsw3dheU/qGq82SO6gJht/KTRuJTK5NToFwniOWgh8m+BuJ+L1PcUinPM9DLYs
NZNvk4uQ1S+Qoa5FpnMp+0ACuJdsxiSpna+OCnTf1t9G/QBN+xLLS6Tdqi+Ox78lmtyUE65Rn7V3
H51R2x08HA99C5+Phm3Ig6pPRyKSv5EZcuffCazKPS+XcAKgIl4OvnyGTL69+9hNcMrocPDxANwL
NsI/H+HGZSl0k+NPfbJ3NuqogJ3sDtHVaOY99zuOXd6GtsMxAbbSOkwieycrNy6twAFdLCwb5dJQ
ISZFN0hYKrus/79YPmnH34EhlGPDseQEOsutSzC0kOWvX020au75vb3NboqnEpOM0KBajJdJx/DI
tNO3UpQlh1oFpZMk4/mMD3SXj+GxndlF54UVPbSe6ESVWqrKwAtmVuC3p+8Ro7Jscxi8KOO/2O9r
Yw3o+CnNo/XIKUizjd5ZU0hY9iBN/+FRe4r782aYyWHyA1unr+va8pYe5jaXWO0XpHQbBq9ZbOPh
skXZlBR7zkedsnYVEBxeD8vWtGmcEQ2bGDmcsnjlbILNgocC4aLccoGJGJKjT8vBo0YPeTVtHArP
FMAEcc0Ysb9BIZdpYupZih6BVa9CAr6shYI8P2axRZFNAwogQtD6HK8jRn/opei8Er3X776k8DDK
PZ0XNplK4elfJgPaB7c/1H1WjxO1AXArpulMPkxjHZL5fQNSaj4iTkauSUJSV8IXG9hqjd4BaKZt
wsLWuQcgX50FOMyjOApWFmLppVmX617I9xHob1QoRbBISr8ppMfagr3+DhOw83oQu4XPw6r9xZA5
H2J+ju9Kxs0rjtKnSY0HzG7hLkFMpARHoMjyoHJ91BFjrmRvGQku+4WSYHc5vlSH3EEp7iiWl5VS
PCgVj6NrYH85tL4b7O4ZtUT4NyYSrGZCFpR79K+dRIC2eSvL5vGu/oWDMSeFsr1RMsMGCPu94voK
JI60kA09U5FiaHpkFuw85JwH+0JV/ZFdydLcQOWWbUrkGVN7YfV46tpIzwENJSXnsJFa8HY+UBGT
8acyyA5ajicE5LhRzlE75lXnFqTuWbtLkps7RBuQS/KIyYR97P3wrufj06aT769w+/h+7PN5Jb0D
R+lgxWYQpSEn05JHQzq+mAyziECw9tPfEby5KodhZ4iz3TVw22/el+ZzKXJEycrLIZLefPcd15gH
+60aR3NkL+6nPkGx83EFVtCRgQc2LPOiDenQwAHq48cgwf0Zm8MAcZbHuRjg3ROSkAupMiMnlRCb
m6kP6sL7c6fzP+QpyfWfbGMaF0fyqh8pr+4uP13iioPjbmeFGwyeQ/IckuGTwyFfyslPmG8Iy9Nt
UIYr6FIRTCpPIrA6D4GCjtcY2BAsSpVk5VQKlOeHibH7khfmeXxV7Sto44ccHV4kZFyAJOm828Nf
eVbZMv4j3tGxy5R7MMqsbdMauvXaOuv0AjaSr+PpU7DQaAEYdAv0Xdrz3AazFkUi7QMyQW9A0RSK
c0Ss+JlgyKPrfy6NnKDXOwhbyeVDYzWJMpSmqJoDH0GrPfeg3A0t7r5diHKAneGingse8/ofbgQ+
Wa1MlA9x840jqgenwr3OWdXJDrEQxvsqjhTUjVbkBm8A44A8IcrPm7+JtVGaNyqBSFuIb+RwgJS3
9oYHQ8WG2vdhmEafFiyaUcKaJ3ks+0wa9BaZu2HuGXw+pKMbVH7NRlTZFj/2bweLYVMdb75mmgwx
5gwDtMZU8tXth081j2VqjJXQTt8eL3cOLlwIlpWwfQrwbls+AOvNNEnYA75ocsKqzsScltEN0npB
QJi4zK8Uzmvj8ZlYZTpFJC3JyI3M8xYCXbc1Ere21zFE4z+z7LBr83kw/lciK1+uTipBX8B6FgAO
qZtXzJdBfOeCwS/9J/PVYLMKBEVqltZLfr/zS3Ah0rOCmwEU7eLeFXyskmpUA+3OA5Uwi1yaX9C+
TCUDq4VkalA1YFbAKWnR+76wS2eplAZlJRh4DfMwAJ5qp2FVYkVDKVQ+h5tGC7ytHlurEKzZGkeQ
eZq5aADEnt9A3fSowxbNL7kxHT0ikumfrepskEnY/Xpg15lxaiRSIOZTu7JC73AejUR0VrQj+SVT
1r55Cx3RNISN9JbBPhlx6p6Q5tJFXQEcKwavGwRSsG2eTcZM3C5TsUE1f3vfYXnHTaIFDb+LqrYY
LfGA85b1atUGHKjiI4odQ/EzSH1aZZbqeyldluE1KatMTD+mPVRKu/t5qe2K3t7XYAHUA251dUND
pbioUFEXhzQ3zcj3/S3m8lIZv7KuKvngwRhuvRt0cspIYXCI8bZ+RuCFuhO6U/pw0anmEY2joBeH
qs0oKuFocDcGeS6F5q4GadYKf4KS8Rk0jHwcfWsxLcKLfLBipGmaa19XzZxktkeDrLaxd9s76Av1
rIz11mjXZldBk/om6JMacgtnBxSQZ2AIkusktq2yga5vZcucofy8mzF1jBrxX6gcnnMTLWDdP2Iw
OM9p+bA+P+hvk0ffAe6vAO0I7ZtKkl6zvQFluW7lplccq6KKV+hqLxGHMOLDEiPQcocZSjjK41H/
CrXW647CDs2Ih9CEqnPjwi5cxdfJvdvtvHMT7c+qtdADd3svuTb37uzM5Cp3UNrD3HG70OqRhNvt
OCp1vSoB1KFC3U6EBDAnIwO81F4hcazNebMxZ1Dy9F0NVR8os3J1VQg/lyT5wvscRXsiGPpOAYWO
YEygGmkpcdS/JhzoFXYO0w7V8Am+IWbdQ8XSOEuuZxs9TRbcbKxU0noD5fjaH3z1D7hM/jgQSgvE
2462xSmhFkEF+SFH5UahjLgbJGVTL8DBNAqxkdZt62f8lpPJeLOc2MPnCGEWkwyK24BRhQDB4c4Q
SHboGFk9W8MF255rbEQtCiIiWmc2cE2lq3q15Mc1E1hh36sgHtp9WjS62hdTtPSqFTD/Wt0GFXjI
9EcgGD8yQdpSWIOqw5OpFP/pM9f9zyiYeTpgVEG8h2MHtpIQFkBhgPCte2b8mVm4UGcUfxOB56KN
y88qBVmpNvCj7w7yg/Ahm7NENXqj4hJDm4HNa4zkQ35FysvMg7NQXL8xrazU2ItUnSPGFSPV9VB0
xeo4fdZLE2uxA5yy6EvJ9YgRMb3bhYsFa/1btn/jhsFkSzNKTjS3SOR3riUjCPZIP0L/7tBKI9UY
AuUcMVsMxGzBBInS+hdbCJ7kUVkeriiTpQEmVRXOwvLnOQ1Xdv8CaBj8go0PhkIyaRla5I5pxppa
HfRRvhbWhVn83YmVi56ttMmDZiwwUQ8KbWcxvvVvwehSE2DAEiK+8F1DO4/igzCYpbHx/4IBW1Zc
S8XN6h5zNqPM8gkjcKjmm3IA0aINiEl3rV61KOc3JAVOEDp/gmnm1nLNhpRLpvwM8XTEVfaKGTy6
Cmp39+rhTWj9ihwaYnB+gwlJIhd6pKwuvkhI5X35BDzI13rfg7xwlZ3xqasnWIU83lXJRxpRXCZO
RlWvKIGefwSkHwManWDQ+Lukjpn9OkHNfp+0b13tWc39T6LoNIJ3MprfXFA+D1Eil8PrO1ePjlV7
nOyKw8GFrCqNkwHCf3aCU5Tl+qW19mqJLmvuLU5SFSFuJCC3VoSl+vFd8xUMuPSvE0349rvRe1cS
FslKEJM3iyZWKGb30p4mttpHbupSMPTf+8BrnhVenmPZupEhsc7IRj5uJwUswcLwkOuDPzjDjao5
poEuXZ5CKwG+dUL9tpbdk6yLM9pQ/8+fUFp2CqjLncZnoUqNq1L9/u0DpEpMWMB8ZgTh11NBX+Ys
RBrC8clSBhHM9ZuZw/1SREysQjtWEtwxNb6WQJu3/pYm31zkevhfnKMisGcQfcvJHq1ajgFIE5NK
ZV8jl2drgOW973d5YEHOdRFu2iXKnxNoxNA9NTM6AeicSAM1X2FSxHRgaU9qD2pCFezEUc4vVbKH
bKXkjgrwa+fg1f2XJWfYPxT3Ku5PzfmpHwt2IXywbFhCHE7vpQqLCw/6TiIr5Y6HEclJuKoEA+s0
HsrCcTZ23C5xy+dpIizB74LnAsR3ijx2uVhCvl9imawPI5RzWJjel7Bhm4ffuVO/iQVmCwJUCKja
A5SGGhKVvREwip/GFqUh8GWc69kauQIFQ5D5z0Y6FQ1QIgwfbUojehTfwWfvx/KJAYngMDR+V03I
7bphT1hWoiUwc5/vy4547QhC2euqaxohW0kaCBhkfvgtaVgdJNloumd9h/mjmzMNBj4We737cERx
uidkE1BWQTdViDwguuYMoQ1LQhyqKU4xVpA2yaIyMBlVEeC7lEznK1R6ELD330e9B1d4T2swjZGA
VDpN1IIEJlSOphvSiPngVae9bGphaeKCtt3VEjF0Kd+M8EMF8Jl0TMIpqle9FFjb1TAkMT7R+373
4JyzPj7KCotaOYex9U6Lgayqn/RCvPxqDM6PWLe5ph4926mCm1M672gxLz8UXjqVAWSA25LhdnsV
4wPm+5ia1JThKTDu+Y0yA02A6aSDwLJNaPomi3dDeW+f9QMORN0ljoetIA35+daHK8PPsBfeuTl5
4c0VYM3s0LykMW3zDjG+5Pfc/EUcADIVp5l1uSvLJwVx7aciK3w7hXR96q7u+6utbuqp6IGZz/zf
1aHuqpdUm/e4y2tynsaZZTE8ytZLHTXlRuWt6NN4vrUMlZRYkogyYuI9C47U0eIr1LT2pkEwC1wK
rlM/2XQh5X4punZnWcW2/w7gx96tHv/VeaIibK+Or3PYlOxrqsdj7T61yY9yg0t89WXPk0QQCDE8
0aBS2iJYnnYt9cnh6ouSWEUOu7TqVOx1rUDHossUqD+w4cBcnjYm9SgSIpY9ogscGpKdOH4qpbSU
0Mq1WolJWNXDT7co3PYfSgerp4EawFpzyFMR6igZp82me/ZeAurZc/sKg44tARKJpDxD/jRy2VXG
mh2V5X6MoMkop/2Kc/K3yKRXUd1YzHn7vrc5hzoe5Uf+uCj8oKNZSvx5LDdFqvp2FK593qr0rov6
G72ihRUtJ5HbZugzjTgr+G1mEUUtraJyrwDRmQ/eldJiYY0G5S8Zr2nhGc46HUlt9vxj9czx65r+
qvnNit+jEcUn1q9zvxtcpHno+Zs7BVbpfpnVhqx2YlUMUxBOEPPdstBeKWPSf1kFAADv6F8/+ZY2
CQdts2kwtOvVQE/Eet/IKRcCieF+DAiOxB1tuSeLlqVARPIrL+/SWY4msDvEunqC01hXVNyg3oe4
aBhtO2rnYN3YL5kM6CIUnlezprUv+l5qRlP2OkU0rUOH3J8lVa+Y+xbHTStCe/zKVLyvIDhL0OPk
2/KNF4Lf3DyL55DzuLImmPW+uJkTJNFfFgsHBrz42GaMstgz9C+drDKaUbp+JxT9YDjWy7cTtLJZ
xQd6l2ayTKkWACu1OpG2dRjeWdPInad69PNI3AN58XSmntlscaAlQi3fShKxSK/UfrECqoUDmBDM
1/8QM/8zOUBmO8lFKk/vSRP6UctTdJHZmMocSPJRK+B/CfywnLBHM4dzXswTsb3mtEDffdeDDRTP
IlBqGymXwIeexa1pANgPdSa3Mg8D713G+hlHUKmV8Wh7rUoDX7ggRB5RlHC8ryapMI31wP1GcH7I
Iw0AILNS06WUNceawpHhwi0ErxkODdKBETuBArLprbTdUIR6Ej1TyTlJb1u8XtAte2+g94VpS17U
+DHFc54vEO362eNIXVPAwDGWoOp3QS7y8OoTept841gPJyF1eoDHE3FLKP/kIPoeydiGXXxNqqvb
cgE3ViLRyy2/Jh22rvpP9VkA3sYtQ4K0B9jKNsPEQeeGfHy+CYlKy9kDdyRILd6Gza+Twqe4+ISV
dqJsWWn+s+xUUst6b0qRkTCSuLZcNNez9WaFUOJP5P7B0olteNjk8VzXBqU5F34XMDe8PjxE+j1O
LK4jU+NeGh84ZN7lj8FGVQDhLcQBQ4NtZSQIwnqVPd7eE4hyh47+wntWAcH9o/pgc1yTjloQGZiS
W8s5hurkrNpjn2R6uPosUJZrKC4C4wNX3OcMZ3LuyUw6KJnEs7ZhE2SEdgQ3ql0QR10IpKiZP1fw
dfNCakOGx0HsAN3ZQo0gXo9eEuT7/KSoQatemy+DuMTAKxpL2cvDVab9h/vRpQ12++aP7BYh9m81
JF4Ga7Ob49xDIK+cwTj5FVaipn/1EDyRkE6nLf9l0Ix8/PQ9l4tIlIBANlJUbrcUvAcD0iNwejOE
CE2JrFDNhw4d6Y4iTlyyB91WhkQ0IgykgXTvbSgEYUqDNqt5Bzf7Ssn2OqT7EvW8R3nxqGupj8EE
DwU4e+rOKgO8OhoI8FDB46ryVTZWoUjn4EOqkVmpATWV56p0uY/dNvw3utoE/vPMZdBAxHQpLQLI
CK8yScZtRoTzQFmDSB6k9fp+0C7Noa85t9Il4R0c9sS+8Y65xS0xE8LE0Xgci5GUAptEltUYTLKC
zutbEJG3vlchcU3kIkT3xAYgW+Jm1FIsR/CXyNLknccAcgr/JsbEw9oAcWXRrl6GVhSowlNxwcm6
OgCxdG0KbRqFnFxrZfIckctwFBUohEYfVfy5X50KXPRlPkBNxFmdu0SRZ5Y4kwDWOv4QQEW/3N5+
7NC7lWpm2NzlYo9Pd7xmkoSk7hVcCQQj6qx662twwPc/0zZlMviQonGwmML9fbugmImxMz/j9iYO
t+XC2KQag6n6tGevZ9jVetqmNEkICzxrwLWEbDPKs2fSr9oBgzJoiZQmx3kX/bhSWdXqXdrU5n48
mvdFVeNs/Zu+2exBvdnBS9RSHfTKOBOqeBqzowrvg/Vgdh1SAk6ZEkNlm6kG3F0LiRiZTW5MhQ2M
oQaRwtVyrwqCt6EFZJarTjmFWmqOcTdwodUksovWbr9BkIc4p3nCRlfPz6TNVW6Yu9U9ws6vBmod
bLhgakWMittbbzhOo6MNkwLcWU2JTki5s5ZSD/AT3B3tFFi1uhtHsS6jY8DUdr21xUybO0lvyrkM
eOU2uwT1ZvEzOFvZo+g5I4uVPPcrj9uMkJdjWcR1XRUR1grw0MM2URxzvtr+zJQQQi9w6F/vdCnn
epftGHRJwSuaez+QqVtBEEtP9Baq5Nd755FcSwTt7HpvBLHRcCz6TIpmICBqfVsd50/00v5cVk1y
MZnzgGzhh7FDY0JsJ4k9r3cDPOn/S2i5Nb3PEYL2oQP7uD4r77CBW6VlJaZHPBWjcZKQnawpJk0Z
1Gm/gxrXrlc8OQghLq3t5KemuMqQxxi+Kd/m7WEAbRY0RfWWzut7/wQtVqNdKinzX7QtfW20zR6T
CROPJZMc1yeyNg8M6Pc5h0vNaIjl4TPipnI9OpWVB+7ICCpzoyP8Yi/c9aGpcoQ0Vw/ElbZnbP6x
l+CcumkylbBOanGEECnM+2jyP9H9Bg2iXv6m3dbdZwa6XbDZu816ZvKJPJvR0dBdH2QWvqZB2Y3I
gKBi+jvjHoOq8gbFdc1y/CFHEbT3rNjy2ttmknXuocatO3HFYyor910/nzo+iqYD9wWZMulZeJ4J
Y2EyuQXwxmeAIemS/TYUu+PD7fyjzES9QlpG9drHydUB/rm3vU2ZRHzwUmxBnCgtgyawHDowuweh
TVq+EPQnRiHzQ6+MJEF7jJJ5OxblqsN9jIH3d8FJdBAgBlRZyRaGiZRpJcibpyL2vRqw8qzbrFLn
I7gxwpVzf8nWIDyHCFZy4zwcOYtgMXKJ6aZ0tEtpCVnDZ3BXfjnbBoigrVideOiUn3H6R2aFN8V4
/0FE8qpTvbqWhnP15ssvygeECzxAm3kSSGil/xvTts/tjSIN9hcO2954bg3e0HOH/XjLHR00Wv8s
Ym0+EW2Sy4v8yUjewbKBZHzV3yqCayAYPn7E2GqvVUnesYtV2vtBcw1aI2gpA0NALq7e9c783QKe
xj6FA5OI+f/SYL2l6loFT9nwdfGo84FmmvSF/mc6xeoib1POpDE+euInnNYPSnhZPG2HR3xXh+NS
OoxJtvkg0mqmhOak1pbPF0BYsdJMbAFPL1s0R0JwcbwgnDlT9y5/qwvvYCzkDFUNLTVrw3mPuWVo
YJHRVy2jUHx3KSjlfH/AFh5SHfv+Bjtf2cU9QrNkZQ91gKSBJt+vXZhuA4fm8Q1b4R6QoZDH0o71
sQsC8WSjGZkPt4Va+1Q+9bls3doCGfKREUSAPB/AnHXXWzaniRU7b/WZMErEfSYQyjCHQ50C1gb4
c256VETcO/oJ8WgoNeH739AdZwOpEATsIgJbSTO/bhgXq1ncOFK0KU8XYqjHzM4cRhWrNpeznJ9T
EGcYO1QqXrCdManGUNnCZssCVcEMIegfHfV6sN0dCwuUwc/q952WrLJ3/rflod56YNYT5RVL4N1+
Ov9gOgdLym+fgM1TyhppaUFoeufp5DQffK37aWAbNwJe3Cu3t8Zy2v4tg03epsFk1btrcrkCe8nz
ubHgTGLVQ0rgzwNIslqgH4Ybwr3N1OSgc2HlKk+WIFusnz9+hDhvhthA2NvP9p1PzXsX/Uz0bTOF
/K3YnNhcwOl3BYW5rxsXr+R9ihiCEbboGsJ//7jvnnJ5bkYl+zxqlSHZvGMTY1yFMsOt4msD4Ce2
m+AiIX+Wa3c84pJVnWvZQ7T4ORecjLSb1DrI6XuuIHwYbk6A3n0F6PcNQkqXULG1OToEN6F7tNOF
QuldNjLy7HwZSmyKLBnyYOq6DOWQeVWLZvvltRbTE5ipj4CpwzDe0wKRbhGpfdoSJN3JPKlKpjKj
80NOEJvUOUqv1SDcqXPclUh1F8odnSrzg8WI/evHMDaWHrzgInC7y+q36jYanVIuHJ1uBw8j2mwd
y8dtYrKUisTtLkBcXD2w6bSrretGiQG4nvcv81AeEy10dUxHc8ptRLuIlRHKG87pySKCprmArt6J
wDh340WqoqM5J3r3t7jzZK6w31PivuxEHA82lp/Z9tGhyAZzV88nJLVbcF39jXWMcDBb2mg3e2G7
tQ+rYRQS6YkRkfXc6pvsSBXh5enNugojFOSKNdMCqX+Yg6jZCcqkq8skAlhDkT680HjvufOncK98
uU1uFwmjvzn8q0oyxLiLXtQp5+KH+9HwrqAVLZs2z0N1uUHsPDl1S9SE0NxJ/udqUHMjDcsswlk7
E7nGObzYfFafnbcn1Q4/TTHM6UkTM2W1Ngiw4Grg2TdL6bLw9bskUGK2d3sZT3E+mIIZKViVF7JY
DnwSRSpjsqiw9/8TM3asWLF7++OlpGmoWdx86/D4TcdQLN5x7cDYZicFEBENBaWyKrIU2whxhjLy
Z6SJERPbKql6P+g/cZSoSG0u+G3drZlcGJ1m7AtPoJPfdPEIN0uCEZRbooSwUOlaTT9mMEtJIcMq
LI4PI3thO6MWh0lNbJaSlIz+SoxfGIaxdA4D19RBIu1tvQPE0c32bOvVCSfu6YbDlNHgZOGftxQ6
OsS3slyvGUaGg5yRzTMKjYcvcNU0CLZj2QtnGfAkdnm9aSvepp9fXC2SWQYLBbODNTHvGfcfee4t
gbagh7RrebY/O/g2x0UXubhvim5O9Wz48NrVHYZT9gl87R79eoATVz8vdVB50lKFus23NweKYJUD
ZYA6tjKcqtDUbWCjsa6sDK8gl2HbbyXY+v5V0gMDNVFN25hZKhu27FwubrzOSGJhhEl36Tsh68I5
d+K2gj8+ngYcvCP4QCRGKvohhBYGmbHJ8YVkigitJucqhQ9HX4rCFa+jfqoFPStPEUT11eCR6891
TkzRtysqjr2VAtjLqyAmiblvYykF8PEBdz4cCmoXuEapXIsVyY5Xgv8w9sBBJxDQUi2ot0Un5Yz6
oDuMm/txG7KMXzwZXZudM5zHlJV+v25dKVRa7VsAY/EJ4MYXudSaPqQrW8oPtEVzdF9Z4OLtxuIB
nHeVJeBjyQO3DzdP4dgpj++el82SIba4JjuY+bahQerOhbMhr0P5sZdAo9HzlzJOghyfs/PfJ8ls
elh91VAt1wlgwvh1bHwdFtP3JWNdmLTiyW4xrUsyJ5K6jtAcq/EmIsUbr8AsYNt7gQT97Epdl+RS
qRa/9C2uWAqIk/GtybXa3mh9a9EgQBjo1DT09AD54Gal0MONkw8bCtU2p3qJFKGM/P2fZVWlp6eE
Jfw2V9goi0A+AOD+SbXJPH1kWaeqYiXUrsckq95I0ltkMpeKst9ZUJu36lEsxTsKr5K0MH0KLKG7
ko2XbQummLGbiB6BOoOO2IJKk/5ALFQVXvRPYzxll+jiac2WY8rMvOAjxB3YAnRIGvdObygeFLj0
Z1KQzMKBOvqd2zCljH6yYZiUAg6wZvzNX8njKMiVO841zkRqVGm5qJOHb3FnGvmfKisE9DJwyt1w
eD4wYe9MLPJoPShPxWWXzEmXWQDbcRntX8v1AnRlNLo7jTOkevRkmOCOndfH43Yl6quAdZglFTcG
wA7xrPILIWxEmdL8+uctIf7qVRLBxgrZ+jr2EEcXkhl1pnXkxEr4xeyrjfNbrhSCjToBk0Tfj4JV
G0QeYYO7N/nPOtfk92Yao714NXY8ys9PqJkn4xMSFZyDust2RF9WnCBkn2M2rqOB9HSZEVg50zZT
+9AkzEHK2r5EmXgnC2qvV2JhG9BYYDjm8Q88HGfg9Yf/1v/yLf40x6szuS+613ST8Q0fNW+ReQws
GccLrlmSwmNOKE+3iOrIDPSMjyK2WjBiI9KZvoNy/9VyNUbbazDqwvtSBzqwZ/ZJUCh6wT6PC+YH
1PAtoIt/GnDlh2hwXCs/+BqVtZvgtq54Ckxsc3fXVe/aD42B/bqQG5a33QhcRFpAP+HAA1WWRIuz
UD5IG4d/qIZ6sbGSUKqhJiWH2w5Q0w6uV468NSFWOerF9kOvuukwk+V4ccy24qHuylJhlA410gg4
D9wW0N1Uc9N4yFiyVnqwOGiDM6L/Jy2Mlcq4BP+I2KYSKktu8BOimujNvyIi+XIRe/N1vFiMPhck
0kxuAOzevxt5MYF4hRGoL2/I9pkeVDawEy+ERyde2IiO2zQrJHoGJoE9zhVRwiammV+te/46ZGEK
qY6roeNsi31XnBBA2EwqGCN6aBjj7zsJ7hy5DFZSTrBhaHtIEis48cQ3aLYuEh0TDryVhsSPRkap
a7V0ahcmD6JQJKKRwhXCp5bXDNGkkjyGaa+jMRI8wpOXCPNcnNC2SxStdeW6jyqumZR0d+Zqb7pp
tyzFMaJkkxWyeSjCKmgRH17oNH+s2nZhiEsskVf1JnBC+JqX49wXuAl/ExrqVBPotv0U6BmXbZK1
Lfa3DpOqBStJuiVc0vu9Ha0V/GL7Olk4y+vtK1PhA/DgrSlwSTh51rn65SDE5STDvlddQCY+SG92
Qbc1XKy3CcY6DprXsyDrsDgYzCxj7l+ICOzElOCvPf6Q1WSNTcncjlNlYI0wpB7DygpNjygLZR+V
TAedS6NonoESHQ/j+xztaPA6TtpKxhtPCZa0NlCVNFmAWQgRvnJBseQxZy+FAgreeGzgk+aNRlkt
IOGOByEYmZIoJyeCQmfx29iubOv+kyNONiU5PHbQrYKS6u4vTdlZ0ACycxbW4ZCODL9R+QU+7jVh
soSrubTbioBlbNeXBVrm0q6Twmn2hoenjqMK5TbziGspHwCL/vp3DytM4Wx1eunI9QnexnAcqqyj
Sve37jzKUJMK27g55maer5RQ+H8KGTWGq0C+KQU9NLC93cz4RpzN1ZHVcV1tLrQNOWqYHiZCxt30
w7NwhMYVKFmrind/OlO0bNUlJSG0hyglZDFL/HVUfWWopirsEteofKG+c2CFrCIrxK2LnoovizC2
JdzSS+JmTox/QNt4HDsg0mvVNmskNOHsv+N0JXpHVKKcYgDJh2LYaTGApo4YpRox6x0FNWT+C8UL
AIYUyP6WL4sG3LQwS4t7ngutsG8rLVayioMnbRQ2SnekCXQRCVRrErifYlFft56BnqTAfpvUl8so
vSbM6puG5uYNSJDx110nAgKvQKZP0H2njLD8fAwI0PGL663jVCOvboPsh+sGeIzF36fPQPEqK+Bf
dV/WanzCV/AYfCYS7Sy9WUvO7qQHA33EWwO+pW9OsVOuZ6U0Ksk5mC4W/hBWG3i7HVkGx6y5CP1O
USflO9TY0ce/DPo1TyeRvVNGXzCHcnGMyzJ6b2djYxShuK5mLmeXYKAiaPA1TpZQrQ+lMph2JUJR
ecM0CGJNbmji7onCFz/teqgp+RU3eLIVM9nPFKtcXVNTzP/LliZWenMX8wjdnkSopB4mtgleKx9d
uSqxxxphuiEh1ebvVWZhPrP8trT981dKt/FFT1xFRRNR+fJk+e4AUI+UQ4QjmCS8IZVZoyCkPqTQ
IthPDr/oWIG6Aw7rbjAj5j8ga+dx3NffWUdpxHHoCWQJ/wKcYH4JufljdWnD4lBUboVX9MiPtp/v
TeKqobs3yGKDYKeJmDFKiKVh1aZPWzRSuijeH5PBr7AerQDkPXt0Lk85DS8MCFy8aEBFNfFmM6hF
PI6RokUYUsXXYOlkBoULcsm0a/dLdMf5Y3Kt02bn/YvHnNwjeZPXohLE/t7aFrMyGLqwNRl2xi19
mahkTNcZHdc9hhx7mIjmWlZkb+hRVxgYh8xoUkoMsT4kZcc1jQSNfEuSFNPUuYmqsE65B7QiAJFI
De6Kgn7z7S854VHhO93qKwcyjWLpS94/b9NB5xFChcIV8R9oWlvrKKW800rTIxs/GmlBvWYzbBYg
S+wSkC55KwI91Iqh089vyW3+ZcvbG8RbahyC0ciOP7gjkXCl9d3ek1pDBWAI0n3EUyYWx6PFBheW
iU9QnbzFO83IWgEYF6sS/RdBwSXTT5jsmkurx1AQjXGVrjGlZJJkxVz7bJYnJ10JQX0BszEehk3J
JPJwP4y/VD25ftbzLbCtsXWhNQ5/XtzEpqGHaOFoaBeYgmC9EZ4wJnf/8P0DhdANLj0fAgovIBA5
cJW1BfGsmJG+krNtdZc4Pf7gyqJ3koh180nMyVRXv1hO092FVE+jYzq5r2GHba/Voc3p0XmlVzut
dhSsfAWfYLoF+0K7tCqy1bqUksIHKsOcf4rJBfhllrjLnl6hTIJIr4ptDJ7vGbgUUmhsfP54PUUl
amYq049IZ3Q9Ac8jF03OJciOtLBcJhv6xGxHDPl77Tl2LKQa0iwOE4w9xHYDhOQ4pMUzahHnISMi
8i3us8hbtaJ4VE7lH1y0rLl9SYailg1aHHQ8YqEplZMUk3MhKgUaS36rKX7G4GbR3aZ+EEx+wy5x
L39OYE0IyBcCJ2kAW2moRVBVFQ3t2giIf89RzpCaAaFQX0OQnfbjLNVdFdQl4qrDBICTm/7l9FRr
XmMaLwCe/C5DmX0W44VqIWiMYKTL7sobd4vSWxpkL0unn8WuKPZd0HjxHfu2sgh+9Ny3Bvcg29jV
h4HgFvg0a2Ll0JhGJJNsmnz9XoO3gOH/ELGNclnyhsDDsBHTwI2OQDxGomkDMKaE1Z4L3igHQTUP
IjBZAYxhL8OZWlzsDWrzRSAj/fTuZoFnTR8Mo+qS4wQZOE4aBdPGGnfKpCrXXYpj/SUjn/7x5OQK
LFXSH20OX6pZEFRJtrS2u05BNZU6onFEyD5s5hLmMUYtofE13T7b3+J90Dk2lFaPUjeenkkU8H3a
6KE4MaCBiKW6rq64kqf17UQsGKWVwr0Y31YeSRMPB2XMCLC055mOqtrRXavF8BCfagOGMhfOYjNV
XKDhWnhCTHX2Yq+A4u7arJzMa9aBDFGbYSGkeyGtaHXLTVTndIBQEHE980wf9tk3cl4kc8VBSKvB
sL1kU6GtzLAp1e4LZRMT1D9SY+D8NRdN2k/n92XIFnqqU+nXNc50ExJ62IaD7rAxfGwVMlXYlFEy
DC2idHx7H9xSeVipDKx3pHhD6xP4AuGxznMaAn8yIPn/JVvZU9YhchASbnxasvrooGsUiLJE/sD6
Q+LYAEg9X+zbZ46/oMXJ+67it5uOZ+BPEzGgGrF6bHezox8TWVRl5ipEuZYUN7gF2l9IPdCF+uMc
QjDmHBxPmC2HMEHGOcS2pyoaETRxMjrZixo0iyN/+U8f0S1tEFsxODs9Xl2cvjRnlb1UD5Bqx6Aj
IXpZk84ZPwaH8n+y6G+sykrVAiELRCpWs3WK22DW0tw6J73uxLg9Ov3b9tGFNx8sM+zTJT8dSnCl
pbkwltqxPk5MWcJ7GjVFs9mM4S+j+U36LyY1Aq54M18oj2/O1u0gPvVTRv3mwcj7dAPdFNiZiQUH
XzQB22wgB3zk7m2GbbeaFuKQ7m99aXFP5DI0F/aR9gjAQdJRAbVyPmPR0HfEWDpHGHQ6WxB0RcBX
oZJ0SBQi7GzcaEQBJ6UHUjTRtEpCJQaFSK6/kIETvKmEXav57qkGBSfZJKgs3T4JgVW4C9fpqymV
tKubVNJH6v3xl7t06Bzm0uyIu8jb8rTCxS1gwWJYW1wlV+/KVaXhUNiScx3VO6Eq4e2Va50tLnaS
1VYv0ZXGD3afc8tTXf2hlU755Cc60EQGVXUCrazKGypu8RxvIZ441P2SuSngLYn2D8NCAgO+aECG
szaZvjTX1BzMhAPn9RDCcYUL/4b92+gM+dmbizMwWwVObH3UFHkxDKz2WlaxBzSjnmBVqOzeY0t/
+V7tNKP/OiyszVcXXwoxi6yRZooqakaMwA4+QDfOXmXs9Cg4WZuvyYi4kKWeWDY8KOo1+7KH5CzU
i/+TQoKljqvEjpKFRDEAKQAfkKgGA9qkyn5IvGOsd784YzaNp9w+EA19NNhSycbXNu/8xW4ZvGoj
h/4SDjWm8ttFfQ42TrAgYopnWLOJH1K6RqRVGevhOoUuphoUKEFGtoYdPGoHw5eUtxt8Jt/HegjX
EfGL9Y9i2+AlVIDug6KceeDKrIFomlLKLCBSquwnr/17NpXED4I5xybqNx8VyRfT9gsu3aYjsSyR
zMcO+dGGZfXNulCH1q1v5htoZzWeX5BEE6cX50R4QBb6dafVeMr0vhiD5kuoa85tLUit4M7MTAoN
fM28W7zIwh/ZlBYG+da+WS5vRohhLu7uTQo/Mf3VqgKCa5osAsrHwyzleZUPws7Z7kJoDeR7unQr
fgTxPB1EEZ0GygP9LoTyGOJfMff2VV0C0lN0ob0jRu+BIbkhN0qvQJYm8KPXLCGqJILF77KoO+Ys
+KaAg2/nC+oBKLKrmHeUtxFYEEUENbVK+VeeC8tHyT40TL7nfyl27dZ3HMpToCEDlPDVOWOWpHYN
JM6+HULZ82cc8FSh7mIW4ooCqBix30yEuZa/vFp/a+GFLqvU17Pj0c73o2Me4EsKfoSygl/VH41n
JCoyluSv0glRY9HHGBmLLJ81ZrEoz6TQu8/sASlEAbN9wFhCx3sQi9OqrvEcNCDt0VKwxUTLLGDQ
FPctro6oXJNnWzh+TaCkcHKR+M/S8p+uib1baeNlqIUMmVV1AEBIo/rg17NrBxNpMsM+z1IKRm8x
mjqxwnW5pvEpaygCWmP1CdRJos9Hm2KUF0/vSVLCMTCrpTzjLPhHWwUcG/UHoMWdRmVW1E08jal9
pcQUd4k5GH6O4VdvV2TqBYP3sZqxtGxhHkKPF7lkyIzp9H0eZaAq0gnMmdGReGazfoSoap9we2dl
V258iSKyG52HY+LZz5v0FREqvQ2EdzrdaiRPscO8QgIc7p65izmZKKs7uKagQWsYswNlgvjkqY9L
BjaR0H02gk0axzK8RsDJWcK68Q0q3naDQDivP0Kve0m1Zt+VVFXDPB70b3r2vTcLFVDC9L/0ZB/M
Ah+WwsHIpxv+W/dIgg2u1dRsiLdCrDt0XlaZMmjPNfA5uNFMojI6SVb+M7uGC0DV5tMnUyqrfGmK
xdVuBwBkDscOM4uLSuft8mQx6+5M048s5jPMsywX8AtGt+SZ9oGxHKsAkYy8sKbBB6q9kOEWdJJJ
IWVDwbr9kkKQL+McfWe7sZ3k6e8eqJWWIHIQfIreWPJ0z+4LNlmKAgLSHTGTECdGOXHCoF4q/0C/
FgfkjhbCKkIIt4h1LMz4WzVnQtnA/AXCTT8xgI1MiICjM/NJN0g+2i196teqXF+7BFTAhrMdALcY
TacNTsrxFkNfVwWPkKiijrNMGwcJHUsfa3ONX/FMHU7iAN1md3MEV8JchPDHo+zgnPozQPTLw6a5
FoakoY1nw0VWu8Us7RTmC1Z3LmaHoN5/JdxLOwQgWFrxeHmYLK9IYtn1Nz2fO3icgarELVI+Okbd
n+YppNB8/2nHwtBATrr6A+C06lL2FHHt3XVP6+YYZhiHOkrCkdh2BSKI8JbdjZBtBq6TBttv600e
PICKAgQwo++vULpcfAjyhA94kA0Mo0IorkfKtfuqECEaEo4D4LSBq1pbAvh6HOoS5BagbGRWezmQ
l/T8c7Mo/ugxdw4ZpTBTAK2AVWTn+q/OMhmWIjI0vweXeIhLkAQaOLOF6T3lUfWh9q84ypKPAfi2
Fjrw79MEmIbSqFsLfWNNkRk2BwqPuV9u4dMOGhc54ZbShWYUuXypcBwCPWZj/AANQAeILbJMCKJE
t2M7iNZVuaDc1IhgP5/toIii57pTWzRPe/vXb51BTEhS2KG+9PIaxEv+Fmg4lrEcpvXPs2wQcRXj
TSIF8cnYA1UKS8fr49Xfq6VNNC+SqVn990Z76Nh4bG4AI0LXSRr5pGeGvF+d/g+jYlYbOAV20XWl
gb3B40PBB4f6a437Gg2iVg/v3KQZ/y9KuwhzuBr0YIrSb3noFTiL6homma55NDZL/NzKdtB9vDMm
PyU4b0IWYk/YXFLvzHv3yJTgZl2aF6QjqgWjV7OT/nLQLkxZ/eSilSVJ79xTYyk1/ODf9CK+2QyO
uxCVG+ilnI9tlsj7YFMn9Qw9xEQkcg8SebND6j+jmtvHO3RTSpkvrKuPGmRDnbwJVwZq/50lDxYl
uB67dRkYwBSYzQ0hK0eOSkeb+CWIm6LM3dIgXfM0MOWze+GSd+8YbTbCuVdG50hJn9crOwJTRJNP
Hvz6XLUC0GbrSF1SRLFygs5XTUa5NgbClOsepPtQd8Mjj/ESd+cbEvXRWUbf67yuGuEUocPbpUXR
WbBhVkYJMNEcqqth56DpAbEE9XAcA+Vd4iBcp0LekhL7OgUGBQZCs5oKxc7r9kEN6QXVKaath9sr
oK3WwaJ6K+H0DZhtSjlBPMU3qbMUHcAWI2q/XV/GkEqBs+JF8nehTrZR/dgOmo42sEYq4l8nQxLq
gOb5r6p2y/APJCchWJ+qe4mKU8SobWpba3uE7VqRlHXe2/IBJFbxeoyNNslurZezA4qmrXY8sbB+
UjuPChQILkoMZ0w39WD5XvAcEC4WjI4Zc8/3L4IEDOjPfbOY5ZsLgZADtUblpNlj/WCdCQdIySln
wysUmXXsh28gdDm2/y/P2yrcDxInnl0zKmk8U3ZxnetLADCWMUExWevGcFRg5B6I95NQASaYAYQh
3sOxALxwjpwyU20b1ny663AOzHVJal6dvUN+xRo4jNq8tMUUoaZgeY3QJAyPZE9nPs8aU/6PvZ75
E3ja6ywAcnqU6czqdqZB6Mf5NIyFJ0JiHGIQjVppS+XKRn+jhNTV4CNqkTzZi5hviUmNqUfas8PG
b/RGWKwhIIZHPQhJ92/6+nATewrq6joSD9QZVkn1e5PgGhaQ6dgoGF2ehWsiiMICE71jc8erzTO6
lQ+5+BippMOS+NDjyzU5CCIPUAoYyeZ9GwLBwmvzTXg8V1ru35D0HbcAJiwjtL59Tn+CMRq+v8CT
bQkAldiB2Dgcby3ujLdjf4VRM5sVXdfcbKYwZJoFA7kmVstmkiDv3MjKECyO+yB5xUs8TCmG+Dm1
q2F4sBJ9h466+usl2WfnV1kLPmG9K4OG+cP+62vGzPJACA3VAqTog4KARj7BB5Oouabzm7zsK0Tg
Gm1BbuxGvtjIbHi7AN+5xL3z7TmzV1G9ZxyJwq1iNxdz5W2/flGbSxEwdJ1rXfQmMa8xXn9fum2B
WAuConzx2htX9e+ZPk65Hx2qyNYr4i2fma7i/ADxEZLqFI9vFr6yH/gBVIHBJ/Gp4MWxyhHtUtAj
r7blY9PNXAtpGZqDzNPn+KI6ckutf/zLrWFBRpEcRyOs+nl8dPE68Baakm9s7yNuE4d++JrLR8A9
+K4EYxP9LfhrHY0PhDnT97th8PuFKHbZG8Qq1vD3EPMGZBnNoutyLhedIcSRO1fMYhG5GDMU4amU
7TzIWeWT021GWOnE7+heijplXQCWwT29YDQ8peIZloC/N9R3aRcCBzqqBqnzjFLV5AR7qXc/lOQo
g5Mx8EsXi/kcWMdyqofJiFGyX/fDeJG000KGcGFRy4B9DteMvTknYhdllsnVdn6DpO9n8l1N/on3
BythukPqlSbeHsJIV0Xavx+msctMrbPDz8qrozrdDH8B1JzSeKW3bKRRAA+3yuGUztve8na/ScFk
QjCFEdyBjD8sDaKBu3Mnrerho5UnWE4f/bZd3fwL31qAdoMoF3lh7LnUmDCwcHOMPpZSSGkOVN+I
iY9cWFLjML64Jau5909mKCoj0eu/51WouceuH/C2KQrcnxyu0GYS7onBB15i0dG9TN6EnA39LTKA
QLM7ZnOY7ua2/p+t8LILmGKwj3p3oydTwSep/EiyiI8vDXdVSPtmsRGRleyt65o0TuwW5hn5ZLq2
hJ2eAucr6vxdT1Y52xiBHJru8P+bo/drLuYC3tnZXncd3iqL2+P0grzVEUzU8mtFP8uWswy3hAHM
lQ6zIqG72tH8PMYwirtnhpPAp8WgxZHfjq8AgHwF1aduHI8+iR0GdlrwFhiCq+IcDrz7cp/mX1Us
wH157STMGQzl1T7i2QUoS32VSGNH9WedHWF8v1X+GOYlDpkqUtEtL/Qc27tV7KWy72xL+8/cwG+c
yg9NiUGhsTIBLspAE7uY+HzYaVd/9bajYgAIEF03WuHH8YOUJwt3Z+MZjapXulhCp3QlwdsF/OJ8
Gh+/TNh7hXXTweRpZFymsZOfO/JnefKyWz3lottZrMoElP67H98AZZHsA4AWwjo7JBt32D/5q5dj
Zjk24euZ0ogFQE/8vuWlYDoLqOSwQ/FtgDZce9g43DAJXg9wSID7aYTUfwdeKQHhyb93LDwbkk+1
sYF2Evbxh0I+jMEZDqLMdbMKpq8s1Yh/7lUBnvHxwY3y4DZgW4oApJjrakblXFE9JRlxgYYGpT5v
fyo2psyXaJH2L+ks0YhaZJJQRvBfwPJhLzKSGbM5D2UfwBkoUga77Xb7TS3DPMNhbo4EymoD/B8S
I9/42S7JK+CFvHCvIUTkDwJHa2HuQr983fsJsesMHMRoPqhM6EclRflDsiErRETT+WMxHexYSI0W
MdZ2d3quXczYOdjV3HYKRjbJ0CiutwwjKudC1K6ktBxeqjJtVe70vGlpPIvzyfwMZZUFsS7Cax8K
JQDUeR6Qti6qPLqEC0yFyLmYV/IZtuNT16Fw+16tUaKDswRa6rMnZak8svB8Id/8ipRKVszMswOH
V1kZkCyBQTnQGnu8sh8Guz2Lk6r9sACnGlvngOgj+xw0Juu37hn5tIDt5Zs2Hm2tWxtem8AlWqHW
Mxooe/gXG3QBbINlOFVFovpUsF3yIAbH5Vv4BT8ccalawGj6zCgJuorvt3GkXWxosbUjW7zo4alN
z638qAsOBCdFun3ONa8YeOOBqihPpLHVeuCc7QZOuTojPLBB13B54NhHk6itVNwHcDAVGRshYE0y
ByHMElf0I6k5OzJOfV2pyVbxQU0Oy+L8Krr9f30rHLcpjLegpX/kWuenVCc0mDmBATCjzPvDTYoM
bs3DFWv17E6+/hZbWp2/+/5y80clVwPEvR0HBQHXydE0ZUyI4QgSNDprTR5lB/CgTHzKdkOyHQZr
ACHieULaL7F+2jbzwxTG5dSRRCDbnMstxg2Idiypvy67veurP0CI6TXr8+btbyC4Q6tSHymKofla
oL8EcJRR0RuzSDShGZzLwHuaIpEsIuSBl4ZLPH9b1cm+UlmB8vyH0BrHcauIJeacKpQjA0qc9HB5
CuJyEUgzopKZZF1i3I+06861mDuQ4fYSDNlsowZjt1hcdt6qD/dWfnya0N4vr7Svpvw5WxejuVUb
kw3B580Teo7J9FpG0EC7OpGhN9R8nEsBy2K2L4Wl+iCEMseFuHI/ratR/whUvPaYvJVd8yWohP1i
KvvR4tonte5VRbZ+5kCpR6e8+Pz87+9cGcj2AT3fGqhV2cxRpkfe+OTHcwG3WChksJacDWnPTNPv
l55HZLB7Sv66/0CCembGOoawQcvDbHspf64MBfG5m0/U7Av/niI/IkO2kXUS+Vja912+2QXNgosz
Mq145wk3WOWXkMzTHXKrQoHoyh4Fjysx5sH1kotCnRrP/PBEfuiEB+kadK6GqZ1tFIFqR0kDV5W6
s9ahKaW9WBwqpuR447XOvodmLE7CCSEgtjHMm98G29rPifEywsMIHKTsZI9isODpzcJocUYJyh5D
LbQRMpVcq327fa+MDERymp7ONV6YWFhElDZ4t1nSQimA2dDYYSRCsok7FZW95+15Xh+SIzoOkmOh
9yUaIPRcUW0TlbbwQwsScZUzRA/B0/NHsMOa55eqAjCR+46mDd31ucdzI7JxvxMOs6b7de+wazxO
ymUTvtAUvBVyplbhdYH4oTL5uonYh2e7Csy/6QMBVShecBpg4e3x1YglhKUMeRU55vOo1N7Mah8E
w7slWI/AIBKQzFATlTLJtOtRlXuhnZ0dls/fd7uQPgCOQYei+yqtbQAdyRKOo26bl98fZJz0Dzim
RgS0KnMK3km1OcPvri8Lu50N/WLuzr91nJRiaXUYX12nznKLhMKgxZrCNQrTX2FmhPkh8KY/fy6X
vWzJTFOzb7RkuoBWoKSZ5+WLLqAEAI5WC0SwpEuP1dorrr8K0i011ifzs048FiJLhwNsKjZTyoFo
4Hivb+UvIvY8F0Gn5D+nKbHiEr9vT0qilDB75L/28BvRrS9WUYVyOcHUnCPySRja8lwxBgtqpQHt
RIVh6SPpU6NJggFztgwRZcySctpKykB2Mtz4xzmbW9VoW9rNuQi+FQYDfd2/ahEMukMqtZahV93J
zofnhvX2CUUuFzhERDHL/EDu+g7qlo+I1WIkJSVGqVN1LsDO+twjOvtxc9MEMBc3hk7Mykhw4Hg7
VKr6BkmK2mMRwoNyl2VPMs1xB7X1Hpv5ZVjaAwShRL13Af8zmUBz7IIc9CNy/2KG2sVg6bMlvnQw
1BvlBGc+KpSIT3wwrmnFSuM8o+RC0lwzaBQOxFbN3OLuhkE15c70D9XbEJwXipaSVzJFAqLbf+Jq
h5O5Z0BHWkiAhh3GIZ2fgWIvOwyYXAxh2gnF2lSG8Ry3mSxsiCQvBc0kDnePqf2S4Jh6kjWRxYWf
jWMlG8fEtesHrvwwguwVgkVLefuPZOWAKLQxpAZY5gGbCQZOaY8iq7oJtAZDF+YYJfAXYltdRUq9
D/2L4XD/Ko8ik5cQzzD3cdENnkkKLLdzuZKZ6CEb+OapS2xUK015HI1h1COljsvPRJ8WgO0jSqj3
+eA7mW10ielHD6U3HyFoP6pbI7PzdjzvBV88+nMjxh0IPYNhVS0idya1e+hWCMSVAHANPLqpKAF/
CScBvlsvd+176z0uEWLOeqU8SUKMtMpdIpKY3NmgaLhlUWFLYcioPagaiCk6Wsg8yLpvUZ0dH6Vz
Gn3RfaJjqEYeXOrcX/Xg9P2u3A8WQVZVaOABgZ9iAOHmc3VQ1GW3lfZR1mVlBIsM3am3j44sUevU
Jo+KpK0P9ZB5ymk7lQl3SZiIWdY+teR6kbm0jdwS0gl0pxEoFTWX26m/XFSi7O1wudHKAYKEZrCy
J7+TxV8khRSQlMuYN9iJzeQaYNz4gP3EYkFP4H/bhizq7fnWgUPx/M7sdLDEubD+urvwaBq6acsy
gly3LQusqKjpz6tWyvzyKJ/QZ4Ix1WqT8rVIMBEnuEkVsfi8RxPvZybzPHHafKNiSUMidjuYttT0
ocS0pfaWd89NKiaLgR3EseHQYRdQcqbpZbMs4bT6+CwxHmmJnf3s5kC4kww+3jxh2Ddq/m1ryMqA
BO9Hs1HsIFqUbXvn3jKYko0EhyDvzSVlQ2ofActxGDsV9IW8SF+LStwLOWV2ADox47ep9+GVjSZG
W4Y0ES02Y0oUQWRMIrqj3gSlaJROqNadxqMoNsSGkO6TcXIKcIg5J2fly1ef0MoglnTXq5euu2W8
mGZ/admQd8LcLVnk2EWQyWrZ2bpLBsB4VS32yi/5gdFG59XyV8EAYpycH1FORUb5cp4xvKXVlzHH
ad2E1D9YSzx/+lPmzOll+/lcudmU4w7aAr/pchGrxI31LwLfr7zrjVZ+3Js7Vgrj+aFOfvn5H4Y5
eFLBuengbyMnf/WuKv+QXBfarjDWiYBUUKVqM+M0dwVqVdYVZaKheYZcv8n7zzs7dA8deqaHtJOy
2rHV2z+fJP7zLL4KMDrwma+Om6vDbRixQwhXxid9/YhFPEkBiSQHazCpr4drltZ2yBidZGwwx/uG
qWzYBGKthn6u/wVhEeE2VIKPG0niMX9H+2/v6xlUr+z3k7GR7X2iJCBER1UJSzsRmQlbb+DrHaUB
yTWOg/0qV16QfViJu/VZcS0j9lbLC9BEzkufiFZ/f2soUzyAA38TXQO3QAKOHYztgNNYBbUAYngW
PMsN2iT55rrN5x4kdpTghiv+TW2gnj5Co1RrWj0U8YBlg0hXJYSHVAGstgWKEr3TenPtDzGwntzv
7UTNJI7lw9fDfc9x72zLtIjnjgCORBF2r0L2fYdR8GVS51pwacMKUfS5fhJBkZzp00DszyK/9WV9
SAtsf7jpwch7aJahtG2sbkdSM9+FFZkHtSloSCcOUp4jpUYZBJuBY/TQTQ+u1X2x4InbdD26g2bL
QMUBaxtoQ76OPL6/65SSTl7CrTg0b5/l95f506gJUJrojgncqzcVd8/jX+EIp1tPyLKhyxRGlnw+
Hrj4RZNlLymR6//N0J8YDdxWF8U7yKafZsNbPlMSGmrzu/Ssyhv31dJ8mNv5J3f+5P55JEHTXL7W
xvEtE6k5qfaJSjyBl7T8WD39iLbQb9nvakgIirKjDU3Qv05KGxrX43KroCqDR0+j+A/oObWLL7K4
Y9ZBqObAJ1kz7aAXwVln6fwPX9rgMjVn3UMiQcjzTT1HVlaf0uKWkqvgob/0zFAAVzTSpBxQKJWw
une6gsIWO3tG2Km7Mf6I9ePfwqPQc7PodJRlJ0bZh/uwYgpNRKPWpyFR6ocXrTl8yFsolvuVSamy
6ExMlSGM8ekvtxT9maO1fVNIs4YIJF7w37qbU41X2K9wl/EPzeedZP1MJTTIFZgy6eLuXGf5elk6
0l1iEbfcIn1M79Bf7VXX7DASKlpKueaqqChx8ZTCOpUx+xN6NIMXUZkWj5ksSFcLlphPdHkUodOK
Pkw4Z+x3GqKoYa2H9dUjCbRDSYnlMK159pROmZ2L7Tl96wGv7V1d6Wfag1i3x1dVWhcQaWlhDxoq
BIZsxbtZbRMN9bLbYlHRfmNnUVMFIyW3XHen/5HNVcC94I3RBB0aH4DIrM/yMpV6eiXY/dBxyEWM
CKOjqodqtiSvix40VXqee2bT2Mq8BgR9ZPERe0z3y8jruLOPF8gCYV/Od74NrevTYa/d161bIG3v
6iawsbFtaGT4fYsMNsHfRe9qz/MclcoPgWSzIPDE2CUXFmDntGNCHtFhfr6cICf4T5aluwNggzNE
sJ0yTkXguPYXUYap8r+D3YisH/bdlLnylKx4H4s40ykTZPmiz2kLJa3WlHCRFdm5/oTzgJwWsyEW
GIzpMnRly+ZQX4860kA1sZN6OP/HcFtXt93yg6u5qLx+IrdHwumpoMau56yVJbWwB99jq6CZvTHC
W+v0J147flvZPTh3NQTslvrJNEm3Z8j2awHwt9INDy5pFjS9HuxcoHYCtfEtm9C2W4Rq1vR8lEeT
zS1/JIxV2vdTUEiBtxuwsDgh7NaS/iRF7AFiuO1OnSu4P1jZ77dh7UzC71WIS5OP0+vZsv0HNkre
cj15jT/95SqBX3kk/y+tvT/L+FwkbkluqOBR37cfgg1OwMZVAW66fUrDxx/AKAP6zrrCISBupiu3
NuW4WPwpOjCUQClAzWkf1JrSt3kpoZ53FuPS+4SD3CWsfTgTtr/C+uefZQJlDZtHa4bFJgLoi/Bl
plYsamJMC0myEOSGC/6Jeu/hP97Qxidybuz15tVPD7XV03a3A2wVC21ZURyWxi1p6B24Sv8/1oEq
qcxnR8vZoVWkAx1RR57CxZWqd2+blHDHAvycDPMGSiO6vTghzROlHXvkdxwsrLOgSgQRdJVxedFZ
EQqeJF2nvJjSl2GsWx6f26fLVg7XlUlCsxxYsXVJOzmAWfBNtCVkkrqn7uw9dS7hrAIBkHgPR7on
VBKcb3+acmBnjv097AJ8v6CBF5U3IWUDToaJVxUzFYhQfVj8cAwmrtmoMTL+7Dudz3gt+thRGcsV
Hfq+puTf8hF4n5wrz9nS13jS4DUE+42CIv2SSICFjvbef8zhtqePd6K1VzVYLnmYQotIYK1E06YA
ia1HYKE15g6XhM2M/GPhhjpLhnCImKxDcb2GW9bQR35a3mvsm8vQHnzdO1yHCtE7T42vkGHCPN/j
I5t7ku4Awd3h7qhqatMKsKtxYKkndBz6ftR6juNqNLKmLGv11PEgijQNHjkushD7pEfhRuj4M60u
o8mvcyqtXtyVBzEpNSxSv/isGADgXiYSVCusu49ZhFxnT0eTswla7h1SqpFOARoq9D1aGDbupdmi
aaUlqFJBBm77OgxNJWUAKqINX+FNaA+TOfIGwomYJpKiyZHmolfhxZa+ITTHBP9Vi4UXNHS3/Oyh
5dfD3Rzr/anlZCFD8rxDEMAYXwsQac9yOkK+PKpbTSZCGmcopplfC3GD9XP3ZTCK8il9AXwBnin8
Zvnx1SFSJQtAw7F7L6wqvMZc0ajtlKtBweXgIGhGeh3sts4+vGxvlHEU82ZwY5Lhra1Q4aPIKPaP
uos+k80AuFuOqWV0AQgj81PFcbIke+LzYu7r6bssCH5j8h1n1mJKWCdZqbKiHdYk+Exj8rbZN4FB
7eKGRieC0ZDXa2MuLkZA/QC/1ckBhh0RiJ8M9gqHz7fxs9KMaSq4r1b4UAI2cS2+m3LDSJMQ1T1L
o41p2DOHdmbQvNiZbPNii/JaiRI3KBRrXuNV4eM1P8G4RflBt0F69W1yPiEm9y6RL+FHMgJDS887
Q2bMBGxoI2m2IKjqYWUoc1CQCcAiWQtW7izpSeYI895Y9uiDKxVcaDWuCDenxyyBYthyU8B1lekq
dCYtLR+nBawDHSwwoH73yuPrU8SOwfbEg5QiYF9cVIdelt9OhtZg29KuQtIzBPIbtkrpPzOB1SgX
OXCm8aZ6pLcDHG9I6w0Yfg2QjxNOcyc30ryRM99kxy7WCuYhz0eeI33abiFC1yGKDD1ac9jd2Vuz
GDMhBHSe0VBzOouQ70MbMhsTWiqurkxiUij4P1gpUSdpPMfIhsFfAUeqKeGZXYCnTQjcBMpW4VJC
JJhBQNd6vkOmXYq/9Tly+nECOwDzeoNI3JrKJ0y0OTFtfeZbadwvmuIGLjvmYX7gsjQhV3fxB+w0
yTRTsK/UGjxd9CrLr62pgVpUsR6Rqrb5JLUanwnIJX9c+3khN3tPhlQcGo8w9VMU7hmz+p/HuZLJ
gx48m2SXn36OqmsNwED/952Rg6vJXWylw2nKn4HbKOGimuNcgON+3cpR5kXR84cTfWXXMsu15JMP
cx4L+S53VtB65VgwTOGLwsBdnJCKCxUHXxSfCiEp7SdFEqEL0F0URk0ET7hRs8fSW0wskLF0nXCf
sZbl1+28BTZ/w3U44l1R/nkGkIYIEwQcIGuujK5QJUvkioVujf+aiIgCe4uT3ZndAXT5qruVLVl0
hYJ+LFWgoOWinWGF6fhB9WQgBE/plW5yuqLyCoXvL1WtMfHS16wU6x0lgOQiylZqgEfD7vpNvA5L
2e7vZagbR5tjdn1tiMGkrG6peZZ9BkbbvXnMp6WtEaadaEKe123EMYnd2bTLK3xkJ7ROixDIHkqD
DeF7rbo1F2HjP8CzOOqCqbq88XnLrlCSQPLNnvJKfd37hco6QCCLBp+BvFMjKfeG3qdPzC38MX3u
GdlabLQpsEETIR1sLYCR7TzAS1r9t2WaP2wKRVAvotl/Bm9bl1Sj40yad4eTqiMjZrFKTgm5erZZ
fAVuCEqSdqwgzWJCOn+5wY/PXPzkhh2UUommA1WbkJj3ri/BYQwGtvzaVmc8M3Gf6ddzfsq/kRXj
/94ag0RVdo3MyaZRIKzdJXK7NS+F4eI5aCxAV6YbtFjrYu4EHCJjFKliWPcJddd0frx2IkMTNROe
MFbHo8qVSTQc8COzr9OKBecueUnoF6a/B0iOigHsoYE0bh/FlNKoZqBJqZlUsvE5tgSyPOHLsrgJ
cxMVYveVSMEKhoiNRr+4vwk4uA/FwV2+u7l4i14djiR0BihUynnnEo22lWYAc1gEj3r3FiB4161H
GuLSBBGwDyLvNMu0zXRT+J332hwn/Qa4KxUDeHRL6AcKovrtS1M3UALwuGktD1XlRhYYTzkLe+UT
XHfi/PS4cVuDLCjUAvMFCRh4nLmRfsg6prPiwqDesnZw/1a7EdN7NlEfPTB/2OXWByWXRbXbKN88
EuHlOiR1Js0IMu/EXM/zxYicR9Fa2VeNad6GCaVxGpYm3yGy/p7ZfZuP/WniPWfAM1PgNRFo7WpT
rUj1mpdLD8zpUKJq6/wbNk7ya4SYu7VHBoLPOgRSou9L2eY4mpmmca2q3aTRLz543xw0Rm+l8T4p
l22AsGLOl4Lc80sBikn6stKdBS7Oe3dJJxBimunN/cQ6qqXojeQwYav1m8253qC7jQ64ee7J1C9z
ldDzgi10jbNJmypSRNMAjr/VaNJVDGMOUMlQdNofw/g54ehMewSvXG8+leNEyjR6BzwCoPIR3bb9
7f2vaYuN+F+n1OJMBvYJG2gFArAC5hT3QwaEqUFzGdEZSmww7Ctk1qtseBypbeOysuZbnwBKHsv3
t2fUyuFk+lLirAHoHzId2/PQ9cOmcArIJBDJ9RKIx2XxUJlYViAOYe74/ckqlQtwI0RVODlZKZuf
AjymZ4Jqn5ok02YNTevihqsN3hsUr0fV9hlMBSN+GWTvyo6Bv6O8nLVBGzmr4Cg/wVyTXoBQEDnj
CVAX8r/yl9ADyVdvAFIOts690o62NG/kcFfwKvpiXC8SEO27GZzG4N+ns02chdaYQ22C364I3SuH
a1KYrAB/B9P1mjceecx2wMToeLwWdzgXoTrhEYRYJCdFlw5plGRftHkg9+VCUHOd3580lhUuozUm
IxE+Ri48kyFACYUHj7Gb/1FDV7yjnZjPVNJ/fxjzDOQbzjLY642gYP7ikG1QPPuIm0+a3FJhaLjj
OIjSmSIdmDvlZb8w6aTIdlg2zOM2TjDFkWciMilSm+BhSld+gIVbXGikFsvfdiJ25Tew+R1461G5
8Yxc57rbLHq6NHQcGa2b61dfJESs3pvNRL7E/+p2HBJEouTL9rjZS3BBFUgaRz9ZBdx2OMFQBjQG
CSsu3EpCy4gClNljTjXZp0apiCWtc2FPLSKPQYur3GzSI3PIXJVvdiz7EcaZCcKivYDAVurGaEfF
a9qhXLxG4VEmEw74/0I6G88d248YscG8C6noIW5a4mU3prrCd0ArFaVC5kS7rwwcGfQS7i7yZYJD
bJelaZMIvD0EyqekimuQBAwol9qBPT5XYDkkWulQjD347L8kJcJ+3occW66Ds8B/LVxtHNA8zobE
q9YK3XrTIx9mO/NrgaTHmCX7TKjypbjYPLhb91AubYa3iXz9u/7BumWIPubKN9cIA7zfQiMqB25M
IW0ZO326MGabFDrtvIoorJFZzYAw+5G2TPilJpw7Gb8gU5dXKp0kebIYCuAACqieH45JftnpMhLB
ROH4qrwjzRPsji/MdjT4oc0/oefmcRTny2fhRrRd4jTFbtTFcxcox9ebxPvH9Yr1kumuYfEcSNbD
EK9MipH/KtISyAAo957StN7Q7sdyncfM7M3KCyrzjbKS96yjtZrrcLDNZlwNdKYCOHWmghUfIq6b
NJQJ6vH0Ds+O310Fw/PSPYUnWyQXpLWh0roR5jTZAyFfJmxB8MVQX4Iy5P7Oh5kpCpLQ6XMjugug
x6ps2rloN/xJ4unArPbNRPJsrYVyaGEysieXdMWGsGL046yvYb5QSmhBh4JgyJJXstzM6FJCdDOf
ZTqWp9A2FdBQ9a5gNo3Vu0mfgIkNrTwjO+tCJPb/2t1vga2Vw8nGr8kt5a9wwwW6+gElvbs1xWmn
+Ma3geKg+arONf0ahd3y89d5BYxGIYrp9KHCBCpy7FvQGbuIdGOkwyW0XDRHu5lAcCTgTGDqBPiN
UC91xMsE5dM/wqzU4//CTdSebwO5ijAJ22IHsFaD5otDIqO7D9G7qQqXDQ9yR4fja0ljH6/DoULs
sAJMZCESEwm7en5F8BCAcsemCDiHR4TQU2IG3uer33UP6/uKsw4F49awgYr7YFRi9PjNY5d4YQmi
a6VsvAh87G2FKw2jYZpFY9E/JP3+yX2kaIVw/N0oeXH4rcKBunwHo6YoFrvL1rF0XtjC74g1bFmi
hE/dApy5Gj9U3RM9elkHJc7xg6uVfqE//hihrH169b10Mc4KTBADzqlvr6wE+6Llwa05ap/7Hb0h
4uQuCroLB5hW3TFuKRcOl6UjZ4H0gxd2OeoYhIpS9PJemZGwkisuh9xCZTWqwaybH47nC7gudQg/
/QSXoNHufbQQ5UcCOyphrL/yp5EJY8ozSjF/5RMN3tkRltytT9uTf83z/CqaX6AiF6IhoUj1BW0C
xzZqcHsJDfmser7AlP+ZlDFFXhKBvF+LTRa0jfuqDpYJ3ibqYRoIVqQRvHXXbvcf3YCG6djqF6C9
zXcpyIa2PqppFlxz9j8kJ3X45JlPxVOmP8gLp+xpL/6wc3HTTXH3A40MbdFNEw3rRTUlJiN2CsHR
ZFyXHYKe1v4koIpXvjOiAz5Dg0dJ+bw8sYcN+VbMDqdHwiZMNnY3Xg7J6AxS8qGBPaJ7OeA0WR/f
LiIspeYcrqEXk/07PPa2zivgofkYKkFde40HvcSCl2Ua9ZALvT8NqPOOzQxzUvFr7coYaBhIv9zs
gY4wqPZY2zl7YhoYxrDBJZrtycJ2ycLCiC7TKe8u3z8gaUyvqXX8i2K6QCR2g5yLk1YNJ39+/scq
MZkfUo9t3ZWQOb3czfdPeQJFY+2DcH9x608P7LxPBWMg+ILk5SvUbfaCL5zivAgKpO/NGHGuk1VW
1muvZ/HtaIX/6uXqR2V4uIFDr/yPNwejvASYBluoou4NibEcHyG+40JX2VSQHkMovizAwqIjTPmr
Qy0xIfhFFdI6MICuj1Zxwi0d6MYTVpljkBu0Joh+LI2miERf2B7wZ2zlVCxE7xcE9+ZbgzP+nbG2
5Ozwmk2Cz3lMhgHPlCPFQ6oxelSxkdIHlI46ZzOpQcj+QJPbf2bc2ZJ24408ldGv0irp6KVPpAvr
xiY37dyXOTFqFAKPWabcKib8AMiuIUzCX4MN074fYsMRSGY37gx+G9MLwWGrwsFotvUzrxLh05X7
gBj6qGqOpHn4FAjwJJKt+ULx7KTLjw6dOTQ0Yzz4lrT1IZ3gq61DxHtFg7ocBZLAV6xKbw/82Tg8
nU+EeAmw4JJuizdwqgO9sjSwgcl4WL7rnwma4oUmVMrDFQU7w7i6fSQXNT1B5AmMOgbsUCfm6YsM
qtOhWn8eJteFl5EDuk+a9U8Y371jb6l/D05+i+WzhDmhgJ/eidp9WAZezcub8VSugNGa09Qrsncq
haKMIw7pYn4hhQQUc7nKr6iATsFEWsiHB24HJr28J7prNRTFgYeD8r9chpKLFMt1NWpcgnGOskxg
456tKW2Vit5obibIoP2hokPW3VtgXxNBxiiaPotscTUusgqd7nNnHuy4MdHzMVFbnR1CD5Yoh+9N
OOJVGH4AMXvDOhuSo4phsnXf2vn2X0m1YykKTh4cMWikGhQ/Rg5htCHvGBeIeG508mvdRiQzdL/1
q9xpO+XBiXpYsKW8b8OcrhJETUbVOVyafa2Y93MzMHl/LFeEibN4Dyi5BAg6Q7BqGiT6ykLnUIKg
3JjyDmW7j4DxVcqYUZ71a3lC+3Ekp2PzubzhJYdZh2Tvk/taxeOiqeH3kcQoRA83qkEQSBxqntlh
JfrcIgcapwfz8kbjSGXHezrQZzOTZPN02DWuDccg103AqqOO+C7ANLHsE8V+0MKE7EhMVt/bnkVC
hcV6HeGB5ojMf9R74dHfg+/o8K4G8Y4hKe8tgv/qzv29LLzaAc9KdHDnon8lV5hGmW7Men+/gdJJ
hYJ60LtVu3+ewSVHvz3BIH+4J76Fm7nGuwQx1bie33mCta3Y/V7GyLcuXgx5vjigKzzo2JVE14sj
sBbI1bsNkKdp543zHmhK4EqL7TKi57oYOgHZtNfPi6utZhtM54uQxHvkRktk+vyxDFrIlS95B1nW
RqZxOYC1ryhPL1hStY170p6PJZNRAYTBNw78BfC0dkFU6wH/pcuf7xxAsF9xjU9udz6lRAha3RdR
WqCxKwrEDy16/tvLt3MvQT8gKJcpmWya/5weBYf+IOHaLUhK0nfKBJ0L6lj3c8rDL58DxkkABPoG
bZmMGXqY9umjoOuD5zd/PC9wvVnqnZ5QR4JZ1da/qstGsHIWwTEuNh/vNT6XUf+SRVFDtwZ7adAw
MjxjKwOCLICHncoh30Wsl/1XIIXA18KbX8A0QidHVVso0okP1exZJxWdhXUJO9ml8rtGYo//d/Xg
puTKGv1JjLSFmiovnyx6/Cz2veC1eXIBtL5bEAhp8BYbhzlRqqfqqsvSWgJKd02WHE5hPWPjAYNP
Mgc3Vif9sJIzT7uMUTIfHqHFK8p1ApQvzSnBv296ZtzCIS+NIEBpG+gCxlwRPN4/DPz+DOeef9Yh
uGtFTi4w2fPno5bO4jY40VhpFDeKxfZIL2X5NeSY90GrAwVxmQhXfjpnHWbChrIbTHRpdqOjkaAY
yBRXtohkqHuWyH+hryTiDRioSK8sOum1ka1YLt9Gd63Q40xaa2WFRaXlUJvF7bXVUBUhARlxOxUJ
YGfXfZvjERxdsoPkpNPXSLn98I9rO5adZUAWTbmkjXaVet+r+Pq/tVXvjdVK/RsgsZx9317ut2Bd
iKsKNapd6bgXxWAwAxeGn1mYawsjCLIbPgvSDQQtuNfaCrurwMBqrehBcgbrRgCCC9fXyBZFBZjY
1Pd95uKMN2pVHquTSRTx4gr9Y52WRzfnNCeqqZl9KzH8Vy2NYj+Tbid1pRovvSEQFpeoRomF7j3/
G7zh7Z43+ciqLtGDDQNpAyhMO/AnkjD99LBdG2DdWK5BAkvWwMMPvBbC2oauArtc8QxrbRLYkh3c
Tf/lZAQPh395HHCSJdBSCnEnv9aDkwjdMEmfgZqxEE38YWhb2mhqE0Q1yM9WP0Erh5eIZVuWyrO7
9vRWSq0R5PKs8ORIQkjkk6vw4l80U5n+hnLGUgCBQgVlaWtQsR6+C3ziWNQX09QtDTKa/n58LXTQ
fvnHtt1V6qFdlKDzsLZ5xVHVArjAka5G8D/k+Ixr6Lmq4p2r+3YTawBPDiWqDxIIekr37RTs2Yhp
XmmGYdvk99W1viTWs8jUMU24g+iAJlx0HuI6+GBnGFWoIgOAWp0eWwKpIdoX5o6TF+drqhjsnzwi
RuK//s+ab09MSNDpC1beUdMs6RifFsnc0SzoElsho1OsCg8g9zDxCAOUC4HB3Coj2gJ5cDiW2vWw
sOjqzDiHwffG5/zYq1PrA2T9vpw48Y0boc1HwpnfEQRRJiPEwhh3fCyeO8+M9sVoiQjAV075HHaO
Yt8ngOPFhPmTMIy58ZI5JlLmSL417FzgAbPh1rdudpqlqkQrBk5hgKmZCykqv6RrtefsqyOzNCQx
4LkzbXwcJwt3tlvO/982pXozmHTii9MtiSF6wA9Wi3zQnppKW9RDp6d96M516nc8PvnLYwxlft0m
BKSno5r1dGK97+pmcgOczXGbyw89E5UsuQqQ4ydpgJdMdp/1I+8gbNg7Rwpfzeba5IDBmk2bY4aj
kifPnXt+lV+Flo3h4LozPDMpCVMwNSi9Oa3n5G9HkXzy8twRSqzobRfbRzuYh/Jsw2mo7MHfSL4k
oNBi7dSe7nH0iwc3gbUEVROrGMm7GbR59NeQz/+R2AUQlgGIEkABMgrHoT+YM3bPrsuhhnTTwIil
cwQbLlzqNvZyiOekdfsuP2NZhNYDs6eTwe6E2EMrJ41mkojxY8ppVNXPEs0r6cvNUtUZPGtP+InX
mcmxn/bFzbJ/TjVY4D8PVUtWUkwGMwj1/2NrBzXFMV6lPXQEz+n3b4kM2EDxGNe5uvY2uCgEBQYn
kh73YerU/wAKoPmQHQRk4jej/U0Pz/HCsVHFc4kcLm0eoJXh7SlB50O2brb2gCo+pLf6Uy/a2jrf
/x0WvisFzL7vUbzfjwbB0tlZ/8JKzjgco1E2Z24J4qxuwZ+nJaHw60tZgndSTp9QI1/LlvhrPGe7
xri7I2WsEDosTZg5ySbrjTcOSK9jr1v/BeZNo919Co+k6My32IjoAQWAhmtUmvpeFowInn8fMvhM
1g5qzJYKBGTqWxXbqqAt65EXpQWWS9Gpuik9cKa3z0BivsgrJshVjHt+4thxgI4EO0Lz7/LaZD87
5pX90wmWskd5RaCN1ndIJ+pCc+8Q9LR3qOIAXj2AQFcrwCpRyoZV2vQk6wLcZucpHxf9gALLgf1N
poZFFe35vLxK0rnqbwGdJri6qp39b17EMFVABT5oIlXlAqRhxwi8ueWcZ5bhlFyb7G8LD9AEH3AS
8kZ4xPu1YvlW8fVc1Mh/jcq9PNBP/FjkfDEH7SFlUyXmCUtRrLgGNvpEK7aVMHhsAsMh4lWSqXUX
WMGL6qE8jLT8wWEN0Kt1pJEIlW07GrtDa6ZT/Q/X0RWoQJfuyt/a3RJPyeVonGFbq0a+3obXSQca
jq0JTxWVgyMjeXNDAKDU7n4U/O5vlVJTTkbUIKVyYs49uJ9O90QqtQxLjGdDgkOJs15QaVCQuWmi
v88R2CNOxIJieRhop2ATtvZHc2gkfQ+QCl//TqZKg8Ip/QkPIcIn/pe9IwYKKXTEQVbz9fG1t400
ot9SAJW1SCTEHsM5LxMr8cfUUwAHGdZBkEB7jE9+ZiZk9iPU9fWFon+S2LVVSOr+ubGUCES4sv8Z
aMDdRxdVUeoibOhmdLDMhvK3whrmxUBqYCEApye7WbkRb2Lnbhn49iluCEhv7KvI7BI0xK6r5oDt
f0Qh8Ll5cymhelcsq2VMAocVvnACqRVUCxJW+WUl4R2T2hwvU+wbIegqdUCwH/2xzXN+AzsuySGX
z3xlB6zB3F8TQ6eRfsdfiAKD1AXVnsk1J9C7M6eDaWz5XjCAPRWAPIdpRdqXrnOzLW9KmQOx+gcN
JFRGEwdt3o6jzkBuemJZQD9qp29KfYgwK7cnyjH4VsAC+nLO572TMO89DX9A9GZHhWL6IZHywajJ
dX0clhtDFGsWaOIF2E21uCcbalvWaLWeu9aEGrJVKr/fuRUDElyYwlDE3cPW3SqcHdLe0z1uryTZ
jSrrpitZtCd3IxJXMhh8KVZ4vTrfsZizN5sQqhNEbcRf0jBau2x2xI7Ozdv5+WaM3oFqVCuG8TE6
fiJ7CeodbDYO+Hh/L6SJeXBHrcsHHr871ymQBCo1higLkLve4eL1QthhE9NUqdqvSlPrHX5yIdcQ
f1WP8LXh3c4OomrEGT3BWxVo+BQUHTysMawJwFOTCa5IIMVUYm0nhIdiFya7hKo2o9tEsMjgMC6D
h0g0LnbQe92JAYY+PwfvEnJydz+iq9scfFUXKDp1GKcBTiWAaDqkwXjS6qMU1+VMe4l720qk0v5/
yOxGvb7t5Ja3fPPEY/CRYVtyWgzB8eTViGlE1xxJ63rraLfAUl4nxcTQ8p1EA/bdOvvsopWZBxla
4V4ejlMCK/d2CQMBcXNkNOSRKrKAEJA9GPpQ6Z92Ig8Qv9JF8Pti0x/ivxO/u7gXgSzKpD4UH/Or
kP0J+lG7rnbB3Q9sQbqQdPpo8owrONAT3eua66QJHSJnCejCKDV9ZiEjBR76DgHoIa+2GxYPfct6
4aDZ42a3ZyJMUVS9OEsvUuSFTeULXEnFrb8cTrnJyedKHSbtIcroSTVrMECC/FiG1Q9tCu5btpIs
pCB0dnFsZ8JZF+WpPsCxcjt+k7A9Ae84E47vzQyK7iNnex+rcIv3oPP2kDnKwF9fQteZBFlCbDzu
xV7MbgmYcAi/+Ec/x09el1mj1lONhnnfexQ5jFiNbUdggC+ziZNKmHJHxFekNVW2CWRH2dfbfaCH
DnJpwRpeWIMEIY7YLFpsIjFhzSdj3RfojeDTXad1nju1TjhxYYU4kOQxxEpwFnp04z1BnhF1Pc4f
fpBnD1YqmPWJ3taNcOsbg77bsNJiRCsAmffrpbIcyu8sxEvnvMstruXDM9566g8EVkJmm+uZnf2P
9Uizf8WeGxlGyw9A134sMF+0NZGaZpNhqoh9FCU2+k1/9x2CwFcDaRJFyGToVldqTTuLMoVt+BxL
qjJbe52MrWV1ZhrAkTspaDdniMDvdMvHUsLJeLR3//qvv5MWfolo8heMyf2RkM4+R/+Qy0Vbp2hc
LaQcphGQxSzE+RtMJwbKU8mTm04kLs+oYXl3Ur76SerIdcvh9qZdzc7jFQID/wWpxXNW+vRlro+M
KqpAXflgEEjQSa+E8xtWu01WRJv1v6pX7Q3aEDNCe6pVHjhbxZXd5mzbQ2nt0+I20LYmqIGaIaqn
lpxN4NWgRgzh6vs7/anIH6OhUkhD4qZWsXmm8W487fOdMCsEP7SoMiyU0/QFV2vCIADq42zR9SjU
IclrAzCoTUVj3M1Ga73FTCz9qKivsncYXO2yTvjc369ER4c3Q8ABAz2wVamu9H6M2mhPS5S/khBQ
thvGTSDnBAqddwnd8T+Kio+jDE0+rZkw3s557HcFGVY9rWDEoRidbIDI5k9H8+WKDCgABX5ZHPfs
QbTAp9lZ64NTqk6BKSdwJVQs6Niiz1q3Hga/p6JFFvK4LaHgjrLYWTFqpRow88AKcKXUU9EaFtp6
HrEAvf5tFbHi2tMSyzsKp7t2MlzMKH+XRnPT6NtdcnmTUSOMq6Qh/0BVMXPFG+3nIJFc+UjfpeC7
4mmXWpwoE6hiOR8ayuWdsc2O0A9gy8r/fkFMkUltPDDWu1oeyG9h9S8Anpb3p+ybdD2VoRrgGdLn
ttHQJZ1RIkhN5yc1oi/aGzDnCyvL3wTh9ffLQUy77OHmbSGlY/GN7qJWlZNs4E9o+6LQKIGkfJAj
pSKo3LflTroAYSeDYqJSDltw25zOP0M6OG1gt2sgolyjzsr2PN53d5WxjOLLjWmCk3nWpy6vHHhl
quqIyaMeqtgSiQK52hpjiFrr7v1dFUl2+QiF91SI6ZPoGxvjJBTdsVfZqV7Q08Y8urwYq/dUt0QU
tNVlis076whjsn5MbxqbnpJ79uijdtIb21VJOmBCUx9R8i7FN1vHGLKbBlPK7IqpHr0FAebAUv2V
PCPlXfp+mhzhvP5bl4pK06ja5maQUz83aMUoXVUSTwhDCMj2HupeiZiDMh84XiFXKQ/HUKbKaIU5
ix94jrwR3gpq5kLR0LFfLn10lKre+LOyYE6DDtByqs+EbRiaeXtU433QWydbTdZS9Ti3wUifxJ8T
WjaZDLS7YUlIjt4wpthu50KiIaKatTz9lujXAwBD8JMSYnyUMqdfEfAocC00bAqioiNq3/4EUSIN
yQVlWG5qAQAM9s1rrrnquqyhsny5Ru4fOnRGdYv+7+MG4hZifXCgWIZbfw7ZAGggMaRFSbc44tOU
wNaoshqI8vU0ctZ6A2C2FJ3qRdCRDUJ4hv7biA7e5qiswupq7cYnunHRg5HN4vRk8zlLbFNzfDEu
NoCB5STaOY8yXQsQ/nYeaAyaOAY+usjwNQ/u7lYShhDU8o6qj8JF8mG21xELEQGcfcYSm1/756oV
sO+6oQwkGqwIIU5HX55pF20c5X2Kx7oxlMHk/otQlyHG5ciQOa2kEKqQCJ7a4y3b27n6DpZjtmE6
Sh2aYHFyL7p6lTi/aBf/aB2pOh0kBpWK8f+0cXdkh05F22j4+o1U8zCGFHVnzWuhC0/YISdFoZzM
5ZJPtEeNCvQRPILu0iKuGMy6sMAgiuh+XttVMZfnHQ1hMuWeLgUzFzalG5Mx6Rggxfp8/q4ubyXB
Xf12kjxOsVp1fsh1abcoWoV6Q/LBScHzeM2rVI/BIou5sQ9gGkVVr10GquvFl0UBxZFt1pf3lSG5
Gt5tJpDklKzajzkOP//ExBgz+wPCPnVNrnSCSfue5Ia17oAMSOYhkDWKBE18jeaXj7YxfCu6/6ph
WUXX8YfDau4dv6reQ6YFK1GMrTs71YiYEpRW/7iEvC/gz7psBeqKpFhOOQpALoU6gUEDU8Xtuc/s
WaqnTWntnTrA9re+vjCWAEeMzlGdznveGixX2WpwKKyB0gA8VPf7xLUWqw5sZ/78ro5I6rpRa7xX
nIeUxZchJICwkPgMFVYaV3RrQtiAqzOnYvYGhWc5vn6wjmAqeDNk2zvPSsGhltJESEVookjNDqHm
fKZmqrSpIElHG+CmzzH10C2Ml/mBvFeYz12MYOzIbhYlkfJeAUtQXd/ot9GPtoKany8Dz1INIBiZ
dXDK9eTCP7MWJ8XCVzfXU8KIXKNFgfc6jn+F32TNjoFzZFKnZ0Ws1CLJMFCwkaJGjw8d2qd7L0Tx
iKzrfKLCgLrW2hon3BU/QqM/13Tl869ZQ1GtoXPLLrJ9LfYuvp+QkiPFz+0+yGDI94XWKuer+aOk
Itt5zmwCk/zypupsWhvqynoR5lI5cd9Oebryez2D+8A4I7TCuNxL9S6CWdOTs4gr6KIJJxko34DO
beCxHNKCGn9XP2BJ3hghFihD9jAoMpg5JMUlHldcM5En8VLPWVqsc5ToP/q0A+27FD+5JErFU52q
bpuUaONXOZ469FJ8k4pRsFAKcj6RAotngK7xEbNUbMxYZ/jIxBlbv8fWozpf/DPxEk8dviasCZPu
CGGS8sRqWx+aPyRlY4TVE5KIM3PlWbb5++5HoP5x8jK5pW+IwekXhaeZeLstghiwVcBp7tfC63C8
xtmQEoZnO+l8M8FJSYKkgzTreXL4ORzPFaRUSptsch8H8EKsCsBwVZsQaMcsT6iGhSmgXf/kVM9B
hTiJNP1GmgrLe6BI77hIauAJJqptVizA60CF0JElkhV/F6eHH6CQ9jvwUVJJ7rwIVhmSTp/54l+D
+1xNSMCNRXrC9ychVfuRtKkYCLvJtcYZqzGl3X8LGER/VwvoEfzapm7GLyvsDTf6+NlfNn9VbB/1
2B34NnkOUXqco8UmfuRMF/AnppU5bTTfc2SnIAUa/7ImVT3im5HRD2GtD1/g+7fRjUTf9wqckR21
oQa2FThiS5GexQ/qW/Ud5+Hh5rS728tW/vzby+CHR3WvQ+ZG3orCXEIndpdubv/2SANrTeCUwCjF
tQwPxxaSBSS1fkipBFzbNHDmsGEoyXXANm2BfXn9bkcrzuqV9YFZxobxUBgZCOPyXPbmQDkBB96Y
Ud4khpfo4dx0r2tlfI0c4AF7EWF5dbX5B/HP1SGslLdsB9BCIPusUmaLTca+7e0wP0S9wvLwO/mE
CmQ5Dx5hPb7T/nq6w9dlA6RpGFag2MdqfsUKKNr+Ih/CqnJFoNajozE6tgCQNl4UBlkkyAhGJyLB
UPFe0J/mxvQpv2FrhT64uwJy3Uju10SI/+Pnn/ot38zn4UMb+VQOrAuz4ytyXCbmNGTQr+sB0L++
1T/BEernYJh08tcr7EKu2JphNvTcbDzBta+82Fd9rffxPLTHyprV91vSIssim3atmkhNIv3ATQWg
u3AhjCxw+RZBkoyboK3y2xn0i1KIc52J3t45kJfEb96pSJNQN+0E/N9sNEwPZDGqozKOlgmgnX7O
+yXM1r8zlMPKWdgNcREQkPDq4SvyWqUjuYqCCamorYOcfVf7OAuIddNGenJsZXeX8VaFnnj35jqj
E4lryzVcQArwyozcKSeaGPjAOT/R2dQjX4Km5h8Pw+ODT5Iacb4ZIyEu7ZllSnKA9FwZhpPqFZD0
NDgNn+m9a2vfoaDh/sqSSYiNh71kB8kYnsTHBjlGcKvr5qcOMzUwxzT9h3pwBTQWuTcSw+mR41r7
wO+qjJQ+QcDfQOPAiM6sZr5NeqlreOqsqR2UhkDAaWXpJY1liYNj1Kg+tU26fqOUXlL1fe7IoZcV
7D7r776DVg0nJJjVoVNSWSrAvyRbjdw/O8motVwcKLHnhng6yqThjODhGr8EhqX9GlPkxEP5wBNi
jmP86k8Q+i13q1Fp9SVnhkr5shp0FONDCDhUEV8rYF6mAQyyVgmlw38IHv6C67y6sKmE2k4MkX6g
ey8VbN8nzFiwc3al7BmfkAWs8fgUeq/KzCPs9mX/oUcWq1m60GUwujpvQKtL90A8o/DFY7KvdV7y
rvyVVCYA/Yq1NzOzpKo2CQB/5VfQ5J/KRfN9wb5IxUyyGsn5fCVtZl0Xm+hriVcf4WWCOd/PrfOq
7kNJ5og68mUQZyR9Ab2sLgACAdUt33EXzoq2Wr4sfoAYkj2mLXr7cuYQQ4tNAMdbHxtzQvY5KEez
87+gymFUElRDdBRtKZCicw4nOjN9uMiJElWquHCLy5tT5ArqQ/jflkikQcrvVHVn1cQndoX7TIfe
gC/RAnQvq71t+aoTY8M6UcFQ0k2gkPakDF9MFnnC5R7YB8jl3rsiT9IHAGkykaSENztaoh/02KRl
LimCFe10l1sm13rV2tLNItE9CbOUt5fjS41iCN2mFKlfpvw7ivHbDFcuO4flPVqW3qeQCSWaIcOf
DTkfa95Gbt2opwlZKFpOQ3yKJ6YhihNK7tQjAKNikrkAwhciApuzwUO0uHJzTOc6sz5ec4IPD7yj
5u5CWWobgHek0N/74AqNpnIbMxbnErBeMtzhnDy+Q85zTCqHi9QYXNESaUhnfQTADoysMpC18VVW
BHe9SolyGhrg8nnbgtQnEfsfpVC21zsceiJVGuuCQM+Ix15N7mDlozMO338gxWO+0w2cJstdWAJ8
q8n6IsKzExVvnAylkFQyF95QXxSj6SfHYkbjFWwW8LPCPVz6BnWwYAtKK60jp8QZriyijVUOSPId
sAEqe5PtXI7wcWYFvZDfB7VjfNFL575qJ86YdVjiwOFqCTq7YxvPjwtEIoYXiihAHbirltHYj2My
NsLWm4lT8Ocnd9wqqc19f3N8PrbaW4jqKGB7iJEtpKhmWxzsn8KmqhZ+sF3jiVa276d1vKizmo06
Ic418jZtIuAWa1hE2KrzXE3ZG8AAdEymegNTFR9qx5v+CLX5JbSVTP3Zo8qrp5t+cLZBnAcDl+Q7
ns5P/3EANiakCKEsUMdS6QRT4g5q554O15cndRCMYgBNb46NxtAPcbx5YTmsoVrcGTDfQFkYBDEO
lUBJCVnHxpQLqq/125BjIi7HtbS1kIppvO7TG9QZrMofo4+Vsub1GwPpceWvKtBhIs6/Ae5Os2kk
Vrrl5OBvnFtSVAzk/W1YzmHQJi1PcrFsTWHnwTCSEKKqhI4oJqKe4iIgu4dgH4hplmoAFjjewxXQ
K1N6BU5Ak48tCDtGqQPNvKlzAa0LteBHsOn8rnZU9EDXZwUy2bHVXDSO8uE8XtlA9IvYRQtPvfuY
7mC3Fq3JXePtDAsd3cPqkPhehHvzMjyJ2kbFIeT5HQMfv3uzs1pJC2hubrt8SyDeFj0CF4A969bn
KuaAPxxFBX3dSjNmXJz9bXu6e9tu3aDjVzeu99D2r2jb0o21YMixhz9xXEtotQzP3xQ5//Ptr/x/
4zYkfchKQATpaQbBEQuE6Jn3ah5tYGt7Qf9ok5N7BS+sKhZvvpdVc5SkM+7sfkdr6z8hZRjqxGcC
dWfD78wEUJuOq9SorXTaPHlACIO4BgajkP0TM9xeFsHtD2YZdcW0fdMS3BhOioYwG7Ug2dipkDo2
tY6XdZvtyGI368Lf/IfpAFk0GxVHCN/FtHE7eltA6xMa/jPe8vV9u9AlM27gzWjre1jn1oURL7EY
LwBbj/KfuFRL3ps+b2XPUSM6yc0ucGAL3Qs3QopcP+agsbRlgU3OavWk2nhE9W8v86DnaplnzohV
HOpKdqXTTAWltdrihxpyzqseJr0T0KIzYkViCRj8VWKJDxzR4ncqxttWl7ATsYxLcfTvSHco14WF
XdPFroWAd3kvaY2mohIilZQfNOpTXJwv6R6PH9HTCTjNWtVw9fk+ucUU3XCrdzaut3LZdLPHkqLO
3hXRQ9iMbcMP4uDQKf4Qakj8CKxTNxjimE5HgUwAqXphLoP4oICx2iLTfYjy61IE/G70MHCVKkmn
fnAHTZThp1CoHe82cl01tsvreve1vUp6JbleEELsWBVa9WfOZm4mtUeY/EGCscB/c0omCBkpFhnH
6pXUz4xEmSiYobPF9WtKwmT0ZksQvd+7kfbab6fJouZU4qZUkHiPzd0ijFXGWefD62C6f2GJxVJ4
0smj2l4sIN0vZ0KYaIO9uHIWzJ8I1CCvDErTHG5qJeVKDkRFOWzPw6D1F1THADj0KPvi0QCrqWE5
73jigM3S07FZWMnFa7sOIh6vyHb1/d5cMe/9myDixLzAYp3hwUbtDw1q8UAhG49cCXRqC5aVGECt
npat88b4UEAsHK0ymQ3E7a2UjefKuO1vrApOm4FfRquNFf6i34bLe1dNeEdCyJDO1UuJUlQB/h2G
dPK6aV5B3oW2qQx8zYUG9ZJncu9tvZeLzh1OkTYF8kWC0ZIzT+B/vhHXxmrZm2PdO4jpL3I3jO4c
n4ZUhYVfTbtR7J5g4i0QmPnqHs5hGRfWqaHxA4ayGn7RJ+8BnxaVHnqTx3yZ0+zHKTWMHKTqP28L
LPHSd28K5Rw0xPX0FUkk7mDdyoi7E5h2bZ7eIrosoBgnHAMMlGB4TvS1+iFmD0f/NfITxmmDFqnC
VlvBpOf8cPbDP+CzwhIeM83HDnkXPZMQtxtprXh15jl7M/CwDngD3o61OWuhnqm/PoiMLQKEHPSP
HsShjfsMH3DNQjtOzXA2J5v88I7n88nM0n1pQa0Ppa435u1pWmI/3nlKMkWWrfCRoNK2Kfm0ANyU
aeV8VYkj4/ZTESvYRraOTZAPJqgC34v3SHt9B0AG0v6/sQLxcT2soY6yulgzfgQk9QadLN48HL+7
8nthrAgJ0qSHikTctaDqFtSI486Q7JvFa8qt8YcMhl/o6PtQPvpoP9sArbthXht5O0pbod58koUz
SIlYKbGTwJVblMNZtdpM4bFGVXv+9uz8JDc6lBJO4IpyAMUR2uvdInW2ARfYQhw0A36WySoInbV9
HRo2Hu2GsOKYDJOFntjdErIOn/N5tgFKvtuRzJOcK2bFHFxsujmAEcdTjWWd+3yXGYoakFlL4UgH
OANabllOokh2XPxrCcpBj4x/qdbfW8bYTWtmyDRc2ZQiGyB84py1LVajIBoT4C0+Vxc4suwVxN/s
UqtS8CmUjRmJhJkZS9gSX51ERqMxGk3nl2zbOMrmumfRrYl3ovU+OkMR6seyqvSy0pVjffovcw/v
g5HbDfFH5mZloXCARC08HkWQTF0FQDBvuY/Z5aAGdVCxRadDZbYLL7na+HEB9VoHoY2xm4SA9rr1
h6+x3/wvUKkDt0/Rxx79B1YAsvyng9hafvdv01clWfdcmaUBNaGHKIF6SzAeQmbDqq504Q8JzwKm
GEU1rj58HX6J5thNiriGC/zCuzS7ovpywiABhE24BFcCZ3y/fJA8Gg9Jt0XBem4tW/sqmUcu+3U2
ny/ay3JyufuhOXiR7Vpg8HXoQG24eHuSklBrGqUPTJw2XdE1haghRPzczCaV/cYDohynY0q/1uhz
neefPqx0wz7VJsCN/M15c+IGQ5mpRpwHZo2bCH1kL1EnMv5QW6PH9OTfbrGnBbEH3S50cogCL0CQ
1dFOj6q5tXGp8Au0dFuigjCPboVcEg9isL4BvDvhAjEzS8mJ6HIJJPBGGdm1hnQ/v7tE47FpbNUV
f63vlSq1C0LfEYB3YpvoLTRo42kwvVrROPjoas2Jb7I2Wygo2/7WzH9lmnqVZtoe+PoZJ9eLmED3
sHjf+1dRFvSIsTIFBLJoD5omaMl+FhNKdP0wTVORWyA422wiIBD0JrtOvfi8+QGg7XcpAFTQ/+rs
Rqea1qGlRskp4BvoLuGM+f7t2THmglHb2A+eN73TMOb154LFFP5eNGZJkj1ShtkOVv44wkBXjWgK
oZqSFIpWPqH7dMM3JgiRbiQccGiaMBrXTQC26X2oXCbOkjQS44QSfB5dxV9RZ8vsmHFrj9byCRmX
bee+kKa63MxGUSHPd73eTxt9l0PUELOdGrb12H5eanx8XLBTZKY30ZOairIXIvhTBPISpz2t1wVg
AMqw7x/jzwfMhHIUQS+zpe5Z4TdIxsbqFa9wWZOflnJO4kNvaARCCAPQ1j+FA4R2A7QKUfK9WFrC
4cy7r1SJGWVCTYpg5IIcF3MpzxYt54H2XLNUKWrt67WQCp6oWhbJrloNUuLST7GBNnV/4CxgFJ22
d3CwjKChpqagEtZCyZ+Act9X7t1SdTI5RB1KV/drQGvXNX2ub4yDz+hWZXAdAXIL6Zwq11uOpvTI
5i7wJpch1B3+3FegdDX6p2V9hnUN2+v3q1wztD2GMsKGnlbXqfVzrFs3ztUFJIMrXgAOMNMdsfGO
sWjqkzT/i6LEaPtDnr5KAXjX/xfBjrgud7IgpyxlXMSlXx+2UvL+jGqZMU8iryWuLqr9RL2D2b1c
sxDFchwRY8u19L0dcFc9FK95Sppr1bxs4OJqkXQIbKnX8r4vAVsfa+1nz1OCY3DpLeLVOQrMYmkx
WDLb6xH0cIu3TkecCM1IpSMm0HUmrLjJ19DX+XAM8dcup+sj9zQVBTxvLAEWKu3p9abvp//s916+
gnuQvHxS55S9YeyOwx4Iz8QNDndoQyd/fWZLva8JzflkFZD+AG9ZXZA2WeyYPN5ah2CaKlbb7EbH
m5MWa7tnm0Wekr/dia2AcyfRKDiRYhJYrQTUhysZulnAq63bcpZ+LNooPzS2fv4pCOYd5QaZuAy/
diH8ZG3+TSgqS74EMpO9468erOmzbjJF+PEer2K9VUh+C60loemLh69cqL4eqm7anjFSKP8lGBSt
yWP2inMiV+0D9EJDkhd0FPUrOmxTO051c+96ezyt6dMshW/TLWE4fIo8gv7UDUGKA1kzRhxpXsmN
BkYMuG8Zu5LKcdBb9yd4jxoQ4IBHU9p4I5BCWKYeCqtJgpylMKJe5WoVbqLj6Vm+QSAFLHiiNxbh
jrbIKpL0dr9AT70zyPNG/r8bL7AYpsK4axwD07mBedyM9SmMKuNHEJaQqmJwQJ+nr/yfYK1DuOOQ
Ofdm8VCRS5bd7roB+ZLEq5EPBUNM9lBAodHhYWVoo8HwAXrCnNa7Te+QtGZ/A+mzaWkmPtN6zaJk
n3E5Obf/uiM/gVi17/FOgWZGmK9EbujNsrnLXmWcI+X8arYt+vIoqCIpXF7zx9ni2jOmhGoqUk2Z
B9i8jo/5tkeyyThkxU9Q8ALdrefkzlsRe0Ava0VVJ9T6nrK/n9zPuNEWCNBEtPHZP4pQxxKqQF7B
C8BfybrUhxnUi98aH9PMkxyZM7yqBDMl6/WxIrvaP8vZ1xudt/j6ADf2I+SGX6eYxTFZ8eH+8yvh
BJGRXFnaYo645WIhSzUlJ82Q3rDwFDDUMsIclKgS6+fVGc7BpcKZXpl+GM5cV2SVuqEdJsnV1KZZ
FDinaQjPcW/fyUlKZPFBlTFuhr/R7Wxuxv4Wh1UyOZVoMqqdSMlv4MOwGriIrMiVDHyza0BS69re
Nq1cs2iFAE8rJ2Cuzm2+0dAq7TNklSX8NRyg7Xvo3yyOKKSsarViuE5A4uDbHwCrFJE+MMmQ8iAM
yGBywINv7c/FqWQFvGGUvHbVZiFzmkbC2qvui+AlWrLGSkJ5Kd2+rIFlFj5k51ZyLWtElwXUVreW
wVrb13tUj9satUmjuDLvgFZUuTARHUaKCofJgeVx4uNG4kwAFWRU2XWCRN/wYR4XiniOx+Cq8kLn
jpLqZV+34R1YN7TkEGTFW0HHDTGKi8nM29iwxZJB4F9/J840xmRw9cMt4LevYJwbYIoY2lZYeFck
tEAGJpTbhtq5cSs9Jx5IzhbsfxQdJtWrEa+4AgrsojkpqfqFQqaCW8V+NSUipAX8X0sDJimdeGp0
NJa3/ZnyCBxS94IuJ+QsSXdedH/Rn/4Fv0x86LRJ3xWS7awW+TJsW5znMmWpJUlTdCFF4rqFEESH
4VBVVi/DO29Mv6SwGgA7/GoWilqqGyPpFhtyhT4nos9upB8TKfvnRoUn99RwmADfqzuB2DFJ0dsp
mJuT2m1Xy+tsYivmW7DIhTKs5tTzgY4DBPpgLdhwwkyjw46FSVi8XA8xg7biU3tiqfU8geHUVw6e
eT2BaC+CI2SCntFoUrA0Vggndz95bN3XjuqP+NT4IqWGzWcSF/3zuOECgj6GFQ20cwWwstu3BYq8
YvbgRTO0t3lrBaJUtDv31831eKgXVfm0KXLi0naDuxO2xikGoXcnNTWwyILq61SrQW7QrvaOekk6
4EMCOIgqkyTr49MsnfQEs3VSL91BXIdip9s06JHOFGJmZFroKJkaXZBHeSUg6H11CRh63VG4p0XJ
4xLiCyLqVc6blTvCburCWNT9BKSxCsXHhz0hg3p7Q9LWhQL1U2wFOKhMifhM03CXjR2QKfdnroQn
gt3tal4DIoW/ivrMlhQwNwbzQ3fndJlev0cHtEaU56wFm6ZNrhNXaokbtuERgBt/zQ/Tqlmor53z
Ymc4EYQPQY9OolNC+DwZQ+dvFrBHN528YFUfKp99p5hGVkHrz5CK7BbMBhKGjiLHIpVxvy9OdxbZ
6VX7fIQrn8FWyrCNyjmHOQORLFuZyvM01KfVy0pVjmTe2OcaXZd+w4O1RyZQa8sXeBo0oT+T5jIj
X3YwgmzVZAl68GMxv2kC+5xzCcJR1cJmv/QDXWN8uZRh9WuH+K6XFeS2EBrs5i/VVD8DPCan1kAR
L50BQx9F+YWLwhYFebgRMI4rmfJfa592YgOwOI6uR6GF+zkV7b5bRKYnKlv4XKkdA6rgy2pPrvda
E1UxZcioiZKNm2dGw03MjttX12qzjGBTbMgLdXXSuMLK9/iIxX/7IYotnex/2yTzyiKMYxyMJITF
XUPXw4DK9o0i2779B25W0q8heHydei+d0PA0kkXWyX3m/bcH9Se2kHlNg+zftGHRWCrb5P7vtM4g
zS30zyYTVvBBwVLaalYwK2zU5DHppEsGMTYVY55jPJjYUIHgSjh5yWYIVE2LwSqjlDPpvaR9V2X6
jNKYlZGU2i1soQx3YZ++X0nUXARu7b6lWx3dRMW1nD6vYG0Sy2la8mrjbTB0rKcpHoyXK5tA3rrM
HSZugJPRWJn10luory/qwdejPSCInHM7rhcXwLf0b8/DVNTcfxyJwLx6mHwzKW+EJBCGxFKiYDyD
2WjAOzvWp74mJrMZ7Wx5q80/J56fLLijkID0o/qvwpRVMoN3pXXRwQ4KSoZAEB0DardhM90W9KtD
MvHX79zaoAdOnz3a3sX49vFm2DQAh+PoTzAncdurCIVhxHb0R50BIlulPxcTlYhq+pzkuPTVTv2a
gJsyL/czOoQT+lwxPCbX57n55/jcm1EK+Ie9zasg2H9JkGoPeFxYp6ILJu/kKsG+vfh7GzTJlWBg
CzorCGaixOD3zdGP8cPs4NAFCfLgMqcjt8Q127T0qEHtNxH5BZS4XCKf0tZQnmU9ue+KWMJ+Xe5Q
QoxpfjAdsIvxYq62L8LuPg7hqOXarsmB1oJZOkvWDuV+Vm/Qc/K2D6OQyDXkPQHAuOjyLiidp7bK
BDJqh2bnVOMgxbjZ8m/4AysEpMGQfOXPM5mIYCoaT08s9dXs7a4AQmZ0xEAH8v5bmwkcXGQXTbeK
xxFx6RajWU3JeYRE9rmcQqQFZkdMefcpxIoz1DIHVP10AZSAk0WZT/f+B20reN+FQoprVrhdnoC1
vc9TvI36sU4f+4ngNjPOlZmStAnV6zB8NHqXStFN7q24RM9Up1X6gGh5iHCD34Y0SFjYLODFe+rj
7HxTF7neyRLF40K8qfu30oDo4YQo85s+pTGyHp9lhYIuEby1MnB0zEkWbKsUVtRHR2LZ2/My2c2h
NFDSfQp/wt6p6pTnSIZzYEE9pqhbd8c3W3Zror8X3sQ8gpu+J0LZySXITlUWX5fXQHi+mH7PQbKn
l7GaF4pCvDmkd6iOepFII4CtHrOHyWJtswsbnN1jfMUTHm5yV1Yqojbr8tJY1YQJRoVhFoTwnfT2
H2HkyonDmUKwsLuWf11cMkfPtqsZSw+0/an8+DAVP8AsgBdst5KeakRZK0Kl4PqPv7eVy3+H7fKL
qXmQL1ge2rTP6G155ivRT7whGN3yGXAwxHA37vDYtTDRRQUvCXXnQwQWwihoQKqNxRNPRpx4ryut
kPCGU6QsK2rpWcVs/HAxBd3RJuT2NpZhVy4ueBRh6ikwPEPWwzBABRcUN+yFvGWkJ0OF/A9Urarh
YzCxMo90mOaPSC+muLsQLZeE+2PuavSPOgmotp0M/t/+MTjkwAhkS569eOBpTBF6y2qsomCuCP4E
ZlR2BrECARI6nMnLPDvtlcDlusUseooUrH8YNC3yTb4T3ScrpmcdX1SFfoOAM+izhVJs5ajkelDa
JKruBDGNeABlEU6NaSFXVM0WjF9K/Hh06zNQ/4p1/aBqFcQAMw70bI/erOe/DCSUG2rXzHSjCyLr
BwNg0+dydPIBkGynugZ9DYj0+Fb4PorNe0dSQ33zql0uvpZzy3YoSamgNr7yeqMfVDSc70wjdC7Y
uklc3285i+d3AyusJiMAorn6kxYqdHcq5fHs67mrGQ4/c94rRVf4QYSkWfIcqHFyX4cDm8f6uX+1
8lTe3ZbwGLLJVh7k4DIE5G6VtQUVT4ohrC/ur6Vq3TqWk9P3WXAp19GYc/gb5UrgpYgAEdg0hufO
ydN9z1TSC31RWRJd9zUoUyQfEsjkUAL3J88dQZIF/UzJvkwjvxUSfKXiY3jg7e4RU7j5cUgYejex
dCM+k3OMioFGR8YarfkRQ6dOkiVCREOUtJuJGp4GPz2XD3y8geuv+iUJ9Ty0OUshgi+KiTDEtRXO
IkXsM7nr3wMyYmd2wpt4NmXvuxkGlA5tev4wujeMeHIHRexVJere9J9q1wnwtk+VXaMBkBB4fKoC
sGyisCV21APPfQBArnCxXddTq0rlgOlkMV2UUswqvC+j7A8ApD6KTUrZFZONIXvOnxFH6FgS+x4j
ND5TzGEr73c5Y7+o5gBKIMvlvT944TP1qiDtL47fKLUwSTjCw+XIWO8CobXBu6oIW9DiAMYxQVs1
BLQ+54sN+5qYfnQbGzpSuRQWLSwAqjkl/G3u+ZR9+RuTEFtsTDav1d9Q66a+13X2U9GUXl5QxZL3
0XNAQHb0JRzaLGNlNvEzsxWP54OWYgcfrJA3aWy0rRQnYO7kdp9zOtI6QOuKNfKkK6D44xDqXj4A
FOZyTRixhec3y1TUh212N7d3riczyVvNtpx/4j2GDj4lTlK8ZmF1sjHfd8D3sc2Gc6B3Yb1DxmHt
EVPzO6hlo249lviOxVoOCuZ5E5QII5PM/49PSl0ySaLzT1HI3zDmRZYc1TVXcBzywwJD4rx3XwBc
TY/+F3YnT8bRE/WVQ9Gn6s5XQU4MpC6OjK3SF3YeGX2QecHwGn3r0UebZBO2jEs7eWz7miYHfPE5
YMo7ZqWDVxQBXrqQwWbumfPoka1Ny25urA/rwjD5pmQGLKrydJ9naO6aEPXaoJyoBkN/aXXNWX9e
ow74c0bCneW1kK6xAbWeZVDbFm577obt4R+nDc5iVEVBWtfeWI4lCWN1Ok18FSLAfCHp8WdM/rVA
T5io8huHxdjggQOYiJF1U/x6sl61bAOZs1tLY5k6R5cFyLDZQkxU3Gul1DoCB9KcHe20Ku0Rlg4e
BnsGc+2AX1d9IG3EGjbNSZ2RlDldEZGENOjLG3/ve5RCv4HhdFTxaY6BA6CwR6tj74mDKCRpbLri
Rvme/+AraZwHRs9bPMJMliezade0fl4+KyFrkCZN928gGkKDnSfWj9G46DF6CcfYxvWPm8KcHxrX
wfhznW+JBXubCXW+4SxHpgFHdlmkBogeylAtL1aMkLdQ1JB09Ftz6EJapL7qV0Q3z5aHfYpf6ChE
ugNHKkcikTuFbxaHEb5CpWEXfQ/j97EiLDJOVtUdxmVU4qhtuS0+Ze87vcVsBRMXKzQPI+SCzEJS
HHAecj50KlNsT50N21kbMU0arbfaYM3z+KbFwUynoWvAm8s5/dD9lZnLV3TFTeiTuzmlYzOUi1Ig
2L3ZlkzYD7TyTiNUpjVfp15h4RUsWq32BEYXpONFUFpwRxr948evnfpZ8bdTIxkaVe2avXBt/XCl
3m1WjyNKSbMPW8QD2gYim5H25kTCpAPjjXb1ZlzZeyi4WZpmeROkAkKUsvIYHKnMu/wM+RpJddc/
eJKtDjsz/Ksmn2Hw0mzZUbr36VcXg5rDXygzjZxkyIA+Bw2+3wVbK4bfWP+CC6CPtj1+VQsYkymg
AKFAIaEVcNRnbzMtNfMFYHBO/1jO3eR/75a/ObNjkxcpg0zyH0D2n9SAuiRE9l3fTv7q0h6u7FU2
pVMOT9+h+xbRJcMwApsMJZA4cGcFoIy/tbTFGnBZKKwfIA4a0B8IEObS+vtWYdVgPVulb4yMsjWU
ZWxKQwuvjCkRiKg44eMxAKV1opGoAbcC/FQBISmv0VkwDsQ62Minklk7RumOLCO1/2XshEtR8Rdn
r4UQ54ajRZjvjGyESzaaBDnN1b+fXjgINs6uXdlQjgsYAVvkjvda/7AXF6r2yKtjHRmIJMeOwgaX
7GFbRO1xcvk33YrIkUQfkLcQ65ljBIRTM9h2/KR60Lfsa438fzx8EIyLzmeOUtAbGT3iCdztlfM/
zOaxOYnHDLiF9GCCZQa5I5BVT2Kw/zDInhvAexdKcUMJVXL2IO5skErKF36wzmXGdySWQKtUd1ya
+ijjXYSODS4/QoAeB6eHyNaAqBVo9sYNvPluHcEhGzHfWtUzjKGSBYf5Lc8NA70CFpGp4Y4P5B83
rREQTc5PwkNtJPvVQiJhI1U67nXAbd0Um0eL4fUc8cza2iIghSbJAQoh3PxLyiXHeg27YSAVm26f
JrTm/jExXxp4R5bL4efXx/UVxfyqCT8fyl12zpNNwNQvlwVYZ8yQUw3ojhkg2cHbJkcj6WyRztzg
DotC+rmbmqVwdloB1vs506flJ/jvxrQH7fegw/gT6GywHNAWminPtu6nXAAFNUlNl4d8giJpS109
d0hBgXlAuJbL45ATe3CvOP5bLtnMWm0/hzTsn4hXTdcYLStEHq4dZ8sAc+Womz/4LSGft1smxXoI
V9/99RKm2qXXvoQ4FUCGCuXwwVV2J3CIzRmMXfqAhxYr9WrhwsPxKLH9K2dzzwOqOIM7ZGfRMrzT
8vd9qm+ZQBfp+b1jQhZtpCPAJu5N1wMExZKmgU/JuMThL1uYqxrppagzxvGIQl9+bhEDp4qrNnzq
OsJM6ArlpisjkVwNg2oO8rNelqapo7l2Dq6el03fRqHH5nA+8Vja5F7H5mRY3gLiLrItehMAzkwl
h1PPUKmDqKh+26KOQXmZf1K+TZFg646FBQOdtmYze1PgrtLTVJo6v2/UvccKjpl4/4LovWxnpoE0
dXeWKAUlEpVy5gPZqUkVnDCnPcefdf2Gz8p6YGdUJ440a0k50y3anvYRF94MEHy9xiUy1+/57H8s
UGEUNTkEi2L+dqB3aQEnedzbyOhIQLnEmIazKWcGmuzjfvS/h9SFsMP5YumUIjLQPao3FM6XWMfx
n1SvJRIAUl5a3GataU3MlihDCk+CC5aDc5Ovc3YBJuC9gCX9b1PDxWA/VQIupB2caUvTA6DNKAbL
NdowXgb1/Jpht7wCnRadnrP4cZ9RpBB3o0EwsAkAyx3ibzROnqQlQ4CVJXv0gEHYxUgOohTfwmqW
Ws22rl1J8p9GvXxg8LzAX8Ng9PzJ8UT/mKfd/7pmGoLSuEwDRyP7BF2ZDTLPy9MVlaoRrg0uTxPj
/3gdO4nBt0d4MnMxsR1IMFeB2sttk4TUS1Yj1nfb4a600ySbUw4K2cPO3jIPxUCo0v88X419tb7G
oWVpLtuGIDeJfnYvoasEXAFyPAtN55FnpdqyVltcofDPbIc218scjJGTwjaOiMdtahqofiMCCfju
KwC3VqvXmegSOxrIkMt7T5DTw2yoTgCJhuZ2QCsHBbb8Tqu0lP/1gS+KNp8Q2vBwG5S+9B47GcP9
ENxGRGk8f4ohnF3dpWIUxcJJiWIxQMK5X+PLpgtG9kExiMKNS4o6f5ex+o+OqEIg0uCe72WIVTUb
+SVdCvhNfsVTYEx2yAuvzEt1chL1IZF4IMgjJ8fYLPf/pPaSygi5JXckWF4lC/KX3/H01fXmp3Ei
qL5mt5sHSVfcyHM7AVg3MTyVGBsKQnPfVBR7GIPzuJwP6jwccOCKBwaRxAF5u9OrJo8yXkKtigGO
LjiMFnosWomqb4mH2CtQ7sEQPrwlyrmSY+HpavSca1IiXcK0tJVMfh3Bp0G95odRRAIaQZM/YR59
q4TQFwFc9K8Dxd5DubXT1tTY85KkspU6GTNaVgP6yMQ5zjft9Io2Lr4OhxeF9EP+LPpS9pO8vpcW
tB7hhf5s8JWctrRHG+a9G+25me/TSN7KxB9/he98pxNjgVKxFROU0NROMhaWYJTG18IkfLfvCBWP
GY/IUJ4HweehVFbC95qCnbUpH/XaCkbvC+sDlw9RzwCKskj3fYiH3mffNNO7w8OxMlNtM3kOq3N8
rLjPXbNjiZvvuZOF2uRhNQNkfU9zxgu1cW350heW1cEjggclnLz+KBejtnMMCUhQD5lIA52BL2kM
HotGeYow9rq6mDHzMamYVqf+HhMV5dYWdKmo4FbrREBn0tTmyAx/WZwno/F8b9bYVsVTWAjlMuzY
UwENU1S86fBiZREKoIL1YNN5vUjJWGlYbIwnxn2VXicIbx/Z1dme7Cf6eUCHq56H/y6Bjm1mvv1O
mu1j87HCtA55BzrK2p+zHZzFADni56vRmr69qiqA9XypBs2nBB54MaLlRw0jrWBNSUky0VZY65sJ
HTIormg1yT4EVwxo5zcq8lLwPTRbLPZVew/RH51gm/lO9ranc5Gq+U6mAwk87nzsKK/aRlHAhpED
nNv5lip360C2sneLqBWvxvYgG2KKCPw0aB+crlgBGVgRZY1QcpigfZNTe+R96TyZ7y053UVSI0l5
u9FDouKe+8oo6in4sdSToeQq0jVOVJ1GbmMIRrC8DHASqA1Fd5GjwpLfc+NBwgFpBDgoTrOdddOT
CfcpQDZktlzGmnsbz8hAginsE/gHPioMomWuiyQW+yDIUIA/O2mK/zWOnJdBal7Sg29kJ3TB/czR
yNHq3QXzaFB73Y1rYPAalfYip7tMnTEre434u00iLh2w9efWiw6ZGu/5HJwObITnncfVhlNzNQoZ
DmlzQQYGLu7HkjlxThCk3rqlqfuPwmtLMvs2CsqMT1cowsoGv51kn6trh1ygn+8unoUVgpelfE8e
VQdeWOlzi1/cmB+BLlW7tJ1mmmlKazBcRP5oOpwLvYahgLpZXEqgm5mnRKkCFnCIZ5NlUiYjb2QW
ZjNt/Y4dj2ghw1n0FK/8gaqP/K/MzvFTPmQj3NDKhQpJkJwyJffEM7LRA/sL73UgtQ7rBrp5/WnE
9WjNlgrY22UVIkz/NV/k1IenQM3/M/2jt1lG0YFMrx5nnTJ4SRQWrN9HWcM4apJlg9ITKKIEKkZ8
m5i19ShPT4ck0SdlvRWbNaQDLgZZTMp/d9Sbxgn6aehdLpyAd5ycY6K44RzOFB38W2ai1YhSTzuF
Y3P5jKQCES33HQMEG8HekCBTztFk36gZ+uFjje2jxrl6spLWLZ86ghiAZmgIcan3bWrnZKRkA/Qo
K5xb1jIDcd7beF58Akh/skfbzE39e1x4iWMOayP9QovoJm28nHG3Z3kpnNGbT2WwGW8z/eRYQa6c
A2KB5Fy18qyaeA13nQdyaZOk4btMJYP5g5qJixoxLGjQfevLwjaxpJnXwTxBoDt2zPm53VX7/o+7
HEQH86fWxdl04DpXB4Lm2SviShHmj12TNfe+QhJVftQBW6fakH97WQkZRa6nVGoQ/jbUA0EPMB8S
kUd/6k4RW5TNXhcOg8z/9RwS/k+SYS8VG1v05Fy23dVjygc+c/9a5KWfCeYs2ognoLIyHXi+VodF
ly59qo0sJjsk60VW4tTihisZ0fQo++JVLlRqHmKUkQys3t0hjg+xwCwklNu7TRDmCjGJpIQJXsmx
fKE0b+LqP/shzuOZtUw6ubHwPUdTBqyofRfebmRMrriR9L0IuRr78Z2HmWU43cJQumUh8g7GP3Kv
i/S8FLA5AWzmqjNDU0RuVfZ1MHmxEgLmSq7nnCF5qMLX5x9xom4CJhkP3DjfTSU59H2LDW8w8pj2
7D4NAR45DniXX6QGRIw/Mvx3ZYqocFmtlkfxBwpIQ3ppdKE0WrGyAkxHw9GZW3w/GioIPEwV1ZMp
LgSOetLEoWU0t0AkLaNz2Rf4eXy5enUM9SxpC1y1cf7BqB49TUwacLVIb7a+ZC4uW/uM8aIF1SxL
HNEZvRQ5GlpaaqwBKa0oc5Cd+kXeddcqaPwhqeAzcsSbkSwrUkNHxj+4em+61rz2NX5ym1zn5CB5
2ouUtSS1y/IhzEYwOKhssWPjRKZQg7pJeX7IWAYKZ3VylIcqjXTjpYcZj5Xc26d83m4WL6bLIcob
EYhBlpDyapQPYb8Z756t/HogBLQFAkPO3mfv6Mw6TFqX16QksDGMTGf806hogcnrWhJeIDx6D32Q
MmIIXwFAoMzJLdHb5PoBaqia0NWr+O9ecidA1oiBG2sNbSadvA+26Es+J/W7clSHItFOrCYsB9R3
+zdKuM2aC/hfKf8rWXVPRA4qi1xs2OmIRyB2yuPNaoUiOsSGu/8x0/tZ0SF1jtOUMSG6QnKG6d+O
1pZerJLvR+AZKXmomKAazBKf9elhe56L3IbnedLNMci/PFdfAGxnD2wCj9tir3OTGFYGp2of3YOJ
HKOrEPho9kCw9JqGxpmouEhZFdjzgeq84RPtxPR8MLaip49tHWQ4bRG1MnXF/qb+juuwoZr87a7F
xz0UuSZ5NyZLcIKKyLOjSihn0C+ibHICNM7nIg8rQWIB6kpun3+4jh8GcNs6uAwKckH5Xv6BHIz1
4Po0n+i4kXQd1tXyIVxWcZwWTRyQ2ldRDkO6vUt6w1Wyel93SHN5BRIRSx8mhUQfOzfN6fdHOUAO
IF/ilwjVECL/65BRnf1vYnVnxOeeqjJ6ZivqHgAx46UstLfAlWz0IlLhcGWtkwgb4zXtI6qWsJUu
YhR4ifJ0MLqkw6x7BYMzYnZr2byKXvkGogd3ByZMVcfI/QCqYiFNjcKUbIfUa8dPL1fyHOiyaHZj
domf3AZ1en2XCk29HbBEe/aQ3G2vCQgmmbO5NoniT8tRmTi5r4LaaO5d2w91vAp1RYZmyp2nuoh4
Zhc1Luu4GYa7V2YFCS2jVYQ0paKs4McPDZOJq1G3WAwH/mw/1VgImQjwRc/L2k3oxgesacla7dQ3
YfBGGFV3J8oi6dTJRbpzS/Ziz92HTrZ5CDue53GA9nUUXMreCoBwHOsRzRoOiON5F7R6qAUtN0G8
kVHoB0GbfF31k/3p0n/EjwL9g4MvaPs+CeYF0UU3XTwPm3fOI6Zq+mFhZ8L1OJmLMiQW3fgq/vN/
u3qXgi4LYXS21ttDuiH020o2Dw3lDkX4KNuOiz5xbcYLJIXbwMaIAlbsYOWvktBq7/AdovkX8tM1
EkagD78dJFfAPw9Jy9EV4s6BQaLnorCQp73uzAanYfBdeGRCFLdoWF0tUl3F9XIybfTKU0hmUVCy
i3BXHq4pyUB261OVTAGKxjRusVhtlantq0iReJ1GHkiK7mNqc0+pBw3xEa3e63+AD9HHQgy/LwVi
0gL+soY4ym3rEGt84pJ2wkDKGRDbqqrZXSwRNkzB3meOaRhEBLHsZD0H2sCHIRvDHh+GCChiI7vc
/g6euyBAK77sK8Esowv807svw9mPSss3GUDttgPQ8vMA7z3FDpRg0vwu06YCciWAJoAVKPeWxkA4
uxriZfpfATMUeoidcUiErJ02L1Py8ZKAL32+Wo7PafG0n75D+saFaAjwGSBOZfVLlGDk46WafHNa
G27rWNKL6mbLGHB+w0qsjZVjXMHR5ndBYMoNZ5aeJ+exfetf6kfyVPqWDvM2JOt//aw8Q6w3FYPO
UKq6ncT2H/BBat+XWU9JewHX8mLgtkIBp0Rv3ooSFwpF8xQx1cQdtPjJS3pJ4zgJ1M8QrY7LKFJh
dFlsbDBoTKm6NyX3pW4mEuV4stbC0cBJ2tm9HvbkwzkTsv0I1xgMv9+66n3S2q5ANRRZklaA0122
LkrF6cOIkGOAJDWH/CJ9xq72uU6vj++7S6byCpMDNlAS6Iqhg1Di5R8Oj6PUYxjJw0YsMnzrVm/z
1XhvZspZ64g1OyAOSmVvH/BVSBU96w8d+h+3k6j3dVX5t4mqREMdgHSF4tMsLSJnse7nHI+v4/h1
kslF5JyituQA0IPVnBpsUnTpHQc4SOPIvXlkkvH+1EOBT7NeqASp0GTdI1LF+UsuUOQIi6p7InzL
Lio0oziCqB5x61crmwk0U2JIkgjIx7c9SmePeXXKGK0m4Qnm40IzzIofzxk4jOgDj9zqaqiDTYVl
YxqKu8TQDpHeiOb2PsPiqKeGLyUpb4tnOk9oYA11y0cVt8TlMJ1JVUidSL0ghBZKjIgfkMsDNe9j
SQ4s0n4xMJES1jfm84GoKSK3KLRL+FYDFaklUWYaaye6Uc7xgCuVHHfo4WIJrDmW0SP9TKr3KOP3
omknhL0mb/iQfuj4mdt6H8T11GxbxojCS2IqZ91QyevwQvAeD1dmzTUxLsxE1dcjiPCAmyd69FTe
CodPQtOEiJ70Qlb8cEZVdLuBl9R+txtaO7qDZqVFUh3EwMQ3DXkRc9Z2cangX4rEnTzRr6Y942+d
a/qv/QuZcuUmtx+d+8tzas+qLvPatnS7GJ55v8r83KrmmCZJtg88fFizwAlVfKXWS16PKyteCUjq
uo7aDKQ/LcoRq11vU+NcrkckRPLfE2bZGxkQC8B4cfufYTmqJItjqoqeqgtmLSgK75hxmvtJwW4Z
CszYyq0de31rSXd6OZv8moJLgyNBw1y7o1jyjUVuXs08cLgemUn3IV0a2PrkdzmIqNOpQ54l0pG/
lbIlXyOzLXCWEYyo9oIEoq4bV5dWbBM7JpwPVDff19NblvkkAlIXE68EB2bwkA1vdfVk+gbBug7m
cQ92qAzNuJho5K9/3AGt8iTh7ZruKVoRl5WLB4IxWJrKsiqHHKh3h/tWBJQBEDZOPscVYrifl/ok
htvf2Xehbt2u5n2Do0cfiQHoFSblFaxfoz28unUQv4WyTyjenngdI+KPWz81AUHfCo9/fwVzkkjk
C/VK7Ef2PmefeH/whdVzZ52N3p0WRylk+NHFb8R30zpxp4gpjbU3UVIFwyq1qrNhAXSBW1pqv5tX
GAsg55kahiFJdkpT1ybCWYbIovN7rwZlat8faNQyHqQH1hhQjaVSnihk4SZJ+6O/lZ1lErglqCxH
zPeGJ/q+4JXSJ32TXL2C/GvbQJ2WrR2vZdYHyPjcYl/zuB9XkoYlizGQBFjLARR4IZ7UjvsF2teq
Awab7gbNauk18E4aekzA3EEglXODGrpoOoQLAWnLSdzIuq2eKzHvrzls2p0+LF5VEkDTuTUfcv5S
B4bb8EHQHHxg4d1G19s06+orl4o/5pdV4maOzNMdtJ9HHf5mSvzN6krQot6ap9fRvFnU9PmRhoGr
DSxQFzsHnZ45ZckWcAQj2GO3euk5Oqgx5vfPX4nShK2oO4Tz4H25lB1ni5iBiwC6rI6EL2dCfyWK
7N8qOPpFjGhHuCmoCWvhht1Hj/AES8h7icdO9fonIBcpCWhwaMm5LWNfw9Swki+PnaknqO5dOVgc
UlLbJiTi1CTvZbBzjzC4/re9bZZxWzFEbCuC7DelmNKGg4sp+KWY4RH8BgbSBRzj1T6lyuBoFbcH
MlyhKj45iehnkaKunYpYr+7TG4VF75bWf7IktgwmTC4viF+l4G8scIYveybH1Jvug76moyOssfj2
uvL+yEThyVod8bLeljo4dC19p8Q5PaHrMs/w6ssAyqJoJhfIz3iq5e8yvl1qbV4b+9MB47TnBjS2
IUxFNe+CL0ri0kzVW5QnDRrPyiO31BRoNS3KYrlVx0gENZbZKGIBWWHlfD+lDsQkyiXjnH0gj9DJ
aLnnDFNZmp5CH1YlCVKgVmfMh/PP61U1DSbImzclQsHlIYMk+0lkahocjbnehlEEBTfcWxsWTDpH
Z/V3fzBDlc0IhUujPhUY7e2NHLmXZziIhisXksE0ejxEajeiikrFfBIPM8XSxSBY+8h1h7k18SHb
FmyyLWxvd3y7pt7XZyfHuM2bJg1wJrLIGYC4UMGTyeQy628YKVRVTuOZFhhVoOy+TZpnWutQOZkZ
tOyovWRRoPRwwymHXYq0/yRvjS4WUeU0/4HphUcRlnqfaVAZKtyrt9dNVs8i6sbfX1fg5yUfhmTk
W21lsZn8Imw1hEemrE7jqahzlswTcCuCYOGvnPlfgr7k2hdlGDqqqVPUxD1o2FDIsVXN6KQQXxDR
E8i2KFPNKbjq0VKhYEB9XrS58hc4MhzBGc+oCw6SRpGQSwhnDVZdDx5iExwOp+iTOOs8ZH4my1w3
NaQ4wtVrXKPCAmNqKW0+OekW95zbDJRB7eKf+jNo6cAZ0pkJn+X4aq44tipzwsVzbSeumnlFFmFz
QP5Di1FzA7c5a3q2cfIxR79+iCCuldZ5Bo5iCzg+LSf87NUwwa0GxseaX1DpNtB26PXqiZSEZ229
o4VXwIOyvNZ8MJRezFRFbu5xcWLWv68hw7pnCqVyqoyL7emEWZZWu6hnir0ehZh/kLoImUJPPvAL
NxNT0rnitvOYQESaFDZXsnZjX5+owfFrWSRecg/GXE9cLtkzztfAuQNgpucfC9/38HmklZMrXER8
0OtS01g0vAtlShPyu8+JXyeexhj/7ygbWIFp88utqEiEXYakLbCLZhONpcIGWYHE5xU2WyWFn0PW
t6z3C+v0O7pPoQPzv1sIRTHB4uOj/tgEdfGzFHGy9i+StpaRrKoedFq5qDlWKhw+oLOvBe1o5Z6o
GtxzQ5huoTVxdNHUNAk1O2dKXR8NQP9C4UABo+bzIFSTsm5clr62V3CBiPlnOgw0D/qNq5SbA4Wb
L8S/t+ldY/frHTA0kAE/TiSVProhjt1mIRIFZjTcgYxFvpfufvb+ad0O/Ow7hSp4uahn1oXaIQDL
AFL7LPayO7K1IA3ew2pNIG0J1zAYhmo8n4OQ1V3O6bKhrePtJHpiaRGwd4eGbfGHQDCu1uxhoAZe
AhHC3NJj3V/sYabtayJrx69Ci5elm6noYYs5i1WxuxuNV/KN1MoKZJNMo6nMm2pPRB2BteQrBzlD
oduKAxuUIQi3HPEPVizYPaokMAGNLeG2AjW2OSMMAjoGOYyhzMptnMt77/7aGAiz8ZZY7IyIhl+J
pnuIPcNg1sbwgQJ2yYEGoPsPQrLXwivwRql1jZrjKQJ9U0fa3aD998Wmi5qvrH8zXUgV/uhUCwCZ
RJVTHvtCAADyo7ED52kKKdDsHa9EqOL/28ZHV5onrRXs0QQ8e1/WVrHcoi7NSVXJ5XQau85XkAeF
6i1w7HKnIfajio6gND35S8aSBRB/QNuqCiA5VOK4Nqm2sbzf9Hn6phKZ6Is4Anl0HKlQcOQV5z9V
7UzdFVjvGWtH0RnUhUdjX66QeBKe4fkC0s147vlkmxB3XipKXwHwzaThRCPQleyH4cvm4sWg6vNl
NcUxb870KqLmYD4+V+/F98pS6QBjswbCMHn6rgxnN9w1fdraOWpf/NwzL/7OIBNOcNiddAJVoNKd
JlDMSluCOqNNAh52ouTV50xQs+OMMLR8XS+TSVtDD3eOAVQD+PdqelQX4nFy5rfuPu73nuAQ+YEI
SURTw8/AFW6k2pWAkTR/w7DGXsZRY/4+8fhPYWP02cKMkP5XySHW2tNNdMtZjpLMtimVJFOunB4A
X5bEAw+iWjcKSwcUpBIxJgwIX5hJ3vVl3T4xM88OZf+iiWgwBSTd4Z1pnLJjZtTWk3NaL5hbxb6P
OyifQKexpPKXlhrCCtKtTC9GWkz5SG2x6oASYscxraU3G5GBSosBoJqkqjbyss/c+o6SPPlWhjsh
KIm8PHK68kp6XWWWjlVgkzE2I5rSTFf3ap81IGhu0y8ubHxAGr9PadkQgx4hd3XCyd5w3kjM2Vaw
SJ3UXz8tHxxZHrzfkngqj3dhsOfvGUagUetccpzqYyucgaB3WvX1cAJBOyyWXWXBzzPta96Cag1o
1qnjbPOwGxJ1PxnybVmGjOVQuN8yBF5ngR1HVHu7jbbqrEP4LCSD8B1L7FhFG63h7/HfT2ZRw8Mu
MeLX+jiWAWW00hB2VyRXLOlZ0e/GlXrkeH2VdwMojtRbJdFDHNI21q6nrjKeu4+NHPSqzIM3pPr/
XobIzr2Pq70B2W3Ag7x6BNTKH0lu4vT4J6PaEN87mSVS1hKtAIgk5cZrALsnJeEUpKeBXcB190Wh
hCkBJ739NTjTPzpQtyDw1ACn8zD8vddLJbOvMX1LR76Xc+6S6mG42UtVHOr/ooFAyA8qI5yI9fYq
//SCVQeqaN3OSfYsmIs5iTEulepXRomXT7xOP/PgtikvqsAWA2+2lsmI1xUZ0ae4VG/73qDhDwqk
1+U1uzg0h7OHvN35yeSO1kwee3QVpmqJA++A51Br+sRIOmn2sWpkI49YxzlwBBN++aSFijEjyDOz
/9ZccNE6nI1+9jBmPvxyiyh/XFbHVvlUm7w+QlMN9ZqKIc3dhp5lO7X4vrh6u2oe7/ib9m9c5lpY
xtpN+JZykLLX9LuHBrnRAPhcM+ci4iSRw/h4YbqmoWwTDbUjPnqeS4Y3vzBBiVfDR4PlbgMMsdsd
x+FTQQXtkwyLM/zHz6dWHxxwaCG7jPhmL/tRCO8VjQ1nDoCQi4pJU/YgnfVEu+CFcSedq8A0jtgw
oXM/+P2pf7Gr1msikT6AuHQwuhcSnLz4wvKzupdCw16J4YMi6AVbqAIgf31WVTgYTBmS2HgyQQEL
K8ZinqLXchPsEKMSE626zTaKwE2adbnJTdxunJ9zTwxNpeCndFoGm51PdOgwWaybR3dKSan01AzS
hHSwbajOGcA/J0NEZrh9REvWoQomgXwHxONzCvsr3U+BeOKTfQQ5SLw8EV6wWQNVK7Om78esR5b2
zKcMgA+q/i+Shzo7pgmwlazD3hwB7dM1hOBBtnAZX1edZnxeyYuDQgZIoXBrwIovvQ3YC3J5jiqP
+pby/i7FrQNdmAlhOcDexWxdFC1u3i5xzTXL0CUx5UQSeWqkK0/37AES0yeuM7KvR411lxuAOd7b
3PdPfwVXi1XMvxeK+B4/G7EcGcbNx+wXCMWu6DBOxZFMbcl+zvBDPHyzFJ+wps4dKygrdqfAw4+X
VideRsxO6ILQVG9cuh9e+SML6BKzrsgScJMNNN5Te7VGSkTCtFhcWW2LEYzh7TF5LiXQUpQPr+SG
mM41kkMkN3vhiTOLbvD+Tb5yJGsq3zFqQ7UlhMnv53UfpscWWXYYrdjOBh/q1H6cXLyTusFSUO1b
ga06iReDv4CWyPx/8CcuUHvQijxQ92Ghuy0u/4dqSeQ3G2RWve6IUUKZyPHL+W9xn+nha10I+Kph
j1IWiTuTEPZpq77sXvK2P2tQI4l30XxBaPs/MMJXOO6dWP0USYEV0710jEYE0yQJU4Uz7OG2Y8qT
5bpVA6rhCLpfSbbOA6RpnZsS0goM9NE582GTFqZrIt0xfMM/ULu25xQSmhmfNFYbTGOl5mNNhd8V
fEG+yWr165Yw0Vek42HUQDxv+pm3jsQHmMxAhJKmFk7y/7TbnP26pQayq+HxcK21sRT8wT/1dleW
ZPUycuc9gaix0GZdehWPBo7a7/SHAYD5cn9KH4x4QJiB+7MhKlIW/C9kfjxUr3OmTJEFWsge+YBR
SJ6D0bgAAl30mTjlU/VkM1qgWP84TkvALKDVthWBZQuvRql2OrPDhCBxyh8DMkwoAbkXsBtMVAdn
2g8dGGdsdMp86xxeeFjPEGjsX25evyxCx/9E0LSRGkSH2FIvYi9xV0JIC6f8rJ8+cL/NSgCoJStv
xr1BkWMWxTU06BfeQMvt9g4o++gEiHi8kRwjmzMRnSAzTEnECoErODJxyHum3LB488V11fPbggUU
0U8ssj5ZttPyM2qBT0oUskab1eDuCrPam+x6HJk8M+aoOz1aKTjX/YAgZZ/dOX6Taq3vUINYa4il
eyel0BLvbAqUoeR2DLOzjTneoclHDqkGivgU06Q7psh1czHwFwrBk4tk1u3C8VJw4CRZIKQ+xfeM
GgZQU8SKBe8LsR8X74WqKYvMPJ/QZEp32bedIILc/Odrf3tsK13dibBEu6CZfLmJPh8EFxVRaPxZ
QoqMplOjmRTM0VvVSWy5iudLwbzNvCZCoiIti/MQWJzGVnWm8RrZOnRAqfkMDGKriqDk6t/7Izz6
KCSYDeSfFYfUsQ4FjfiBmd5bWeUwMGuGJOMQi/wmrtlH9JCwvGkEkmC6Ar/Z/l7muoQKwmKPITBe
YtuNZ1onlG80xR4PNnv/vo0rNzyvNqMkZCEVWEpHfMOoTBp8tDCVJBIk8H7oOvCYIZAFaEkwjCT8
5hZskaPUnkWqdroX4J1N6QV/XmtVvbD1ORqP72yJHbojYmR7O+TR/oo4mQqAN9lkm9solnWQj0N/
uIc7h+Jtij8JyO9Ir3CCHAD1IcadsKMW5Y829ZTtOsbKS++wPagC6gRHSzP+SJGgsqKk5Sdne+H3
LSld2tBFIIBzNVhRCgsBQhTW70ZYDG4RKGFcHmcaoz/Y7gQfk/IETIeAHk1TwCl4zxhXyzOyff+2
KA+aP41G0Uv7eA2RoQsbNcw6VTeCs//K24JR5qxE6bc/5QmkC90bZwAphLetDh5KxGeWFoYjSalD
jyKLC1y9h7gfUQqRnu78qjq8O0zLERzrX651Ygpw8z19DG7ikthhuD116EuLpc9nEMzuqxS0r2ck
iTUrvJGAr40WsbC9z8evvh7OTAC1vRZcZNM4I/djhWmJ6ZUBdgeM0+S4juMobg/vCmVJFehqqIn/
obXOzhi4eXvF1Pee7/ZjGbHEnIFnb27ArTO/c2Zz1VJ1daeAFbJwYpFsYJMTwjpWnQzxLjnQSKxH
FXxTmAED2zE+a9ZW/P9MSvAdVk4cMAv7WHVc2AnncH6LA081q7bZB6/5lrnq9jPu+DAWtNcdkF3Q
rvvta+VI982bUDrjbdWd99SHtCJYT23Mb08yIze8h5U2BzqeWPJwbh6hvrVwmcd6Q8294EupufnU
Oxzpm6qzleWxgVusSs4pMuygwiDkTn/23TZAyfF+KtGHXtbOHDPXt/GZAlDm1ixhzcWbKbXDKkrE
N/AR7roTFHBtOD/JWLP+OWOJqCZMVU6Phqu2qChOE6pFkZithPG5rLBHoNfkQCjP4Wa5+nvdyQ9c
cXQYMkkG64dIotgq15t6yHaYxVYj1Gm0xrOOzezQg4K/y7RTtOBE8qqGNFOKqS7vkyn3YIMiOmkV
d9RTP+sVo3/u/WpCodkLuCTP/0Nicgpf122bWK5t3a5j6oxgpuPjnvW6hNflAj0szVjnpVNbnNjc
PH8cH7bkU52w1Zv7r4D9I9VkYfOQ7J7OHPX1OS20Z5IIFOWav4u3/BDj0a8q0ZWwmJMHmphuGido
9tMWiNJsOWDJ/3rXvuWMCF6xWXeGTrPnsr77/UmNg30zuRZZibt7EIg3HZiEX9YjH/FrNlg+iVnX
mvhka9v0evSBGy4oB4aqwXxqBKAmMVoeiTi8fcwHM5fNz+kqjD/BDVMjJmKXDq2SbO9Jmdo1cJUS
PvKSLZkL3G6qMOqSDIZ2OiWzJwv+UjmXaSP/7UQpxEqSnY916UgMquzpVFNOR57J7Iw032CjrGjP
5iu/u/nO7aBhy5bwVvkj+OHDseuwavsGTH1fDZsAUvMZuTMS+QJuSH9nYgXifXOpk7tJ5RF47I7O
m19jVynMgoKeNK2nZkxXfxTnDjG/8k4iOqNIHNpYhUSWgbBPk1+tAuXU7pbuGCpzjF4peOYA+tEf
GnvRH00hd3KQobQvcVV5HptwXeqzZLmvV0dZeat6qy9YFcT0rlSiRTSmFGxVHmSkwnzftPTTtxNh
qNtjtaRnGR3lRqZIKyuG+haicQtCHf2OIpXCvO771kUReEn3R9CeTTk0xT2/ntaq5evMODK2HMYs
1ddV8MuFzZFvD61HBKNO5y10aaoel4mvsmec5gD2x2Lsa6J0BTR0udtRukpwH2fsgtSGYOoCNcT3
G7yO137SL0mYi3iiaxcVuDRv0bX5y7mVcs0xuFtapkY70Fp1ZvzvAjtvALKcJ8KojfDCcUZq6oM3
SAekkcKxxaOcxp+4ByrJn1P2nSspllgYRldkI9FCREd9OgnE2+3teMux0KKaUsqlgQphsRXOBixf
AE17qPatT6ACiHaPC/p1MXc8w2l3Ld5ijKtpbDMOgh4kZvjLTGLOznOLmHBWxsxOl9NSacaPd6FY
2+VBek8sh2ujQoTofg9CFgzlvZif+XNRgsRSUI4JcUTmpJdTTpPRQlzBs5DBtMIc7xrjX82xb22I
Kc1AUKkcsi84krG7GZsUIM2ZFLlLAIX5oRQXu+cvt5ns7qjLEELrxD67U9X3jraWhCXjWUHBxStd
WrEY++MEyrMY/tgibPFgo+qpVj7EiuuVbJIBiGN9AYTCPmHq2fGWZ3KUlOY9VbtBElQqAXpC/JJc
XgY/gXbHWS7pO2jR+hwPHOYqhAheSESJecjxJdk4iqIwbO/+8ajWJM7s8c/R6EICQiQjAxtj098C
pN6v8Kb/cM2X8Ww22fkmTT/MWo79v4rc2jR/aGlJGQuh5Gn+blTAiKpPZ7rnepjnOPXvTVOQl3jU
nsCQpc85XsUBu0+NBuq8ZMo8sFyI1V3XEtQwnGqGSmxgFktvylRCmch+e3Xj1WF67q+TohvXWmnE
oWYV2rkUDZsyHF5AjubEtb82qdeumOWzQyZH2Uz5dFOIm7xy8qQ6MEsd3X7/0sirhaqttuMLeqF2
L2P79q5X1SDWzXhT5yobHGhfrXBxLAsFy04gxi+4VJeLDPW/AV2+deN+uTYU0kX4j7/ChAXv+BSD
C5aEElzzc0wkOKv01Z+2rBRW6Xe+rqUOJGU6ZARpYLSBTPJf39yIt8a7HOxbhY/0X7eCxNFfW/fT
GObXgc130dmMm09RKFRwH8K5sh+YYV0k1n6LASBIKENnQMBm2KFUhzMjQkeXxf6eu91OlaFaUTGY
4UnUX4pEWoBRHKzGINLHYsxPdBj/UCVOMMydqGLbKtFlQAhVX8vip2x6lOlRrqlqfxDIcCXS/mg2
EBYHpsuWfst+z1erdyzV98Fu4H/ArKH4ziLGlrH0s0g7+QFeyoBip7b1xrqshotwSmhSqAZFIXaQ
O1WnCVPcE/z99nhcYnveg8068PnqqL2LYE3vEPOYZNSOYDwX4CLLpK8imQKp6MvwofOzQM5M2UC7
+/NCVJDFG3LzEP1a27pkOtlJFpM0Q8COomvFDabsxLBcYiYBSbY4NrMbu7lwJW3xPhQ1CiciMCTO
wQrAzR8dti3HYcex6uiKAg2CQY7I/UUAga8gTSVpyCZITq7leOVii8D9+pS9Bzjke39kcmH1f9I5
vnnr4nqBSSye/pGyVdQHtaxmL2b/ULikfAXfupYpgT4OrO/sr+fB1rwoqje6g0/BE60oszHlhLFS
NECuvmlmJYbNZLouWwsFi5bg8P7IOKigbmcYGzDp9O1lfGJnXgZcmAPE9XY+YaDSBQVW7uD9+8XF
B+46KYCtUywiOCUBW1rlbn7BgqeDPO8CqsyNOnAHQyvZmypFeaEQbREErbIGArLEFNoX2c13Poz4
9Upk0vpnqNQG8+zNhEzWa4DxeLHfIF2yDk913G+DJx26MRqV3AkKbKo21cPjooKzSqa8usY6WazB
FgPXQro9iKjb24pM4cucTL4Q9Sw2ACwETwBtG4TBBmGCAWlS8HMQ+Pg4tnrj/i8OS7zckxm06IVJ
VcBrMZFxfz37a2HhPr56Ba5/vczVwFd7mzSNbhPav9sjOr7LGBWE5Ey8mqjnzhA+tSy5dJORioPS
TGAUsyPO9O+L5aRIZnnYGhnFDaAyWCB93ILmvq05w9Y2kypgopNQWu7Gp/YiGHbpmIDBk9aO4Zom
QrVFsWxlcntE866FX3UBCY5Tq0B/fY0gFgB1qVvjJgU0+86YWgpK4jEvSr65WYo3JkW4Y8cDWnyu
LlgECDZMAb5DYTlhkr7fUgAyw8ACVhIFfJ+0K4k5ei3yvpq2c4w46KmnQ+Ize1ju7IIU+89OKzs0
LpHb7NeEId8+/fDPztbKHKuF7bm71bjihIYBzHi7snIMgOfqUW3JJJK/rcrllsx+V5KnDZiXoZxs
gE6bBmJ31xCn5Cs2wMI03NOJXhRZ0KJ+uftA0JIFnhf6JYwZgfNW46R3T8riT5gaUOygHnwzQCS0
3Mqi/h25/ajCidLVmIZAkWGJyDJMDoSNUTOG20ol8zr3BbqFZFYI6LLmh/jlTCRTUOIU5IheU3qO
AM51zyF8X0uOQDQ4lO7eYFTdgUthth+pQj40W1XTx2ngQNbB0tlUWrbFbpaoPikACCt+mQ1a7aKW
0WoEMOBC96OCTpXrRTijMoNvXKS+fkmkKXVHPabG2cP5HGk9k9tnwrhrXfsHBg7+OXEllZrQkKPB
Ylf1xPUVe7ipw2L2um0IiqkhIdd4lBbReeDsy+HGJZpP5jEjZPbWSRy5r7aBo1+riNbtSk/FcmQ4
QRkRj7oq/o3FNe66TTDomho+JldXyu8lZY8J9Xc8rrTD49Vu+yoK5jGRZ7nLqBwFYMp2gUr/YyTo
xnoFSWkX3PMt3FOLkaW07yCVgW4hv0M6KkstwT92QMNoUob2M47l4tmsVNzefaYA1lSy/Ahto6yU
Q8OwD1zi5od7vBRFgEOih2FCbaGsJcRzCRqhOGx3qF11dM5NRfoJMx/mY3CRDU9PJQ7hl6uj3Afe
/mVYx28bHfhHIqi8+7t4EgiZHs9Yk3kGApNc92WRhZtQbT7t/9jav9gEuGJR0+FYF3XVlnneRhJV
xj1NLeAMwfHbCCvPLwZySyPJvUlSE62SLxYTdrjGK1v4rmyNficL9+TMdzPM5h4194h8kY/LHSjS
KkMjiEFv5GKuVhwQ2ggGJ4hEY3pIHCRuVlxYYJGU2cj8t0SEIHE9frH6k/p7/WTPSTP0vnKEWhha
NhJdbWB0d1pmROm0a4ekYI1CSfBh7IAS45/hb1yC2bSwZ5IiEvSV8ohDfvyR3oUdu4z7tXdY+eFF
JrNKsRARLigyvk2QcAMv0pz11Lexs4vVySauHoRvUgjyHM+IZUYK9CQIFb280amC8V7ri6Q/+t5H
bp3G7UoVUBcJwi7xjVH+5HsYunz4cd9QUKSA3YUh9VFSYbFxRsGYMNstXwMGMdNG5bLlXTi/OfDI
DY+FKE6qH9K85ycP/KHS1oqp0zHh2fTiNQLOG0brZn8oOuyXrM6Ix2f9NBw3svwMTAlamfPdohB4
aF7NOUlqyhSIfbqolJMw7ZtlS6xzd6r0Vopo5nepVtd7KiXXRBot5A5gvjlED1DW+9B0gJIs3SVZ
JEwPqs+jFgd51Piy2LwYADCMYmuQ7dPXEJVahaLKu69lw6YzdAorAaq3MfI4BOr9JC34eoOWZocK
e1xr7mSwSCaAnunaFaTV5dwmjxlOSszbMgnA/OaeCk/i1J6YIZUHHTXoME+XSeO6p6t6PmGdMWNc
+nBWDfi9VHdF+l8vqJxy+/nkgFnDX2iECkSPumWLLeKtZCp/SiA8aLvmXFdvwReEBu1npko+MRBZ
ENekgsKRxuaoTWTj8LSIAgHYTDF5pn0FybeGKMR6aQ5Ti0N1d1IZkmwmDqwoLiWZ1y2ADA1b2eyQ
IVRG8FKH9LpJrqNLaJrfFfhKloZjvlDvgTr06N6EbYX7rPzm5Zgsg9a33ifbJy17hXBoOYPbztCQ
wMNajSQK/F6qFWRsdXCOMBIuGkuaoAJ1oNWVJu2L6GCZe/SNgIapGi2TRT8YJZxm6YmfyyKSvsLJ
76RDas4tKRCe+i5aj7SmLZSXCqurN3beBP4UaY28rLMNnrC7AZ1lpOLzurIL+GxcTHl2aAcr8IbO
FWPEPYsQsE0Lo1ijDkFc/IWTSJ/4IrF3sCDrCMzCWV45r++sxpZknmF/xVzj8Mm9+HVzhTc3NiiO
WoG/ypf2LQPYESfGgjLYdkqcDjpMgxCQ30qYFtXB1c/I5CHqHvd6PToE9is4U1NPKtapQTeZxZ7b
VSVU3j8UnejFYZL8efA373vFlmwcxUSI8VKZ7XJ1T5x5C9wk+/OnMCCtI4q2VEymZkzaOEVNYPJf
RCo656INxSlZCo9r8SoUpKFJBd58CUvSRNZzsCpLSYHB/t5en0H1YNYWB0OBKkr1UAKzKXP8WTdM
DFPsGmfE6wcFvJVQxUAHZDVtmCVQiJYIr2NK9GnzW3Daxqc1tSLzm7z4C2LLW2UqeueJ4AV+tRLc
OZm98Al19b4LoDIQlcrRF5TQt+9GTDnMYDX92zDVoJ8XMaZr4QZkFRzabuBIt4Q5xCieqgLx4BnN
/UZQg4Z1wjQpowWXhAkKOGv/kQn6biQKQmsvd+6mhuorYOiGuRhWBctJvdZ2dmiwDWbXTMdv7gx1
Yk2raAa5aPGiiR+9gMOMq84TZLIWW7sWSo8WLl8agMVU0G/AfXolFLoQyVrNhbh3Xlaaq5hI7UZE
PDy194R+0WCP61KFabt+7MOpXHtM6dwx6bYYrY5O91ahh6pl9yHdJBfmS+aAGFGDVaUYUn0UcxYK
gjopFPdcDNmp0Yxldno6APRIHslKtzYmxSOVUs7oEA5OkNbRrEL4prna6t5G1ZqGIOHf/mvVS8kD
4EqVkpIllYawx+O8ILO8QrXTSUcSIHOBW0CK6H0hs+yh7b7+zf5PhsVTdnnKP77ULbk4JJeIUgMO
YDQOGOUHHYy0fscQoriKuGBZXEOP0ubKHPzAlCzEgEZXcUVDpZM/o4BEpCpIZ1ACR9APoVcQ+Odo
Skd6sY0IfMWIlz9DvUWX+Pa5KH/z0mb2MpcYQrR/nVmRet2MU9mkr5E3RJmNq/cTrR6ZEFdDlzi+
zpaRm+9fIVtgUWpTr1UBKDt3HmqJTE6QXiBfcxeepg6yPcLCFmoOKsr76rzwxVYb5l4O1alD0Cr6
0IKJ1/CDi488W29t0lcfLTPEf0kQrrN+TxpcD3ky8h8f0HdEvesNoUCz4fGnb2OmnHVJ3Dey01lo
wPY46E6g2zkv/UjcICZToRDg2BeAL52owlSHFLcUmswJ3FwhRlqNhsZYvBeyLRPubLq8ZM8iit2E
Gzyu1Qp0JzosAul9vB3glMV8jEpDJRO9gWKoyIJZpLNwb/JvKXy2tkNIgK91ddc3yq649TJSTesj
UW9NCuBCdw3uE/cg+qULH3PUIrCQubHKqVKX/tECaiv8mfCjnabXb3CLPTfNCfSwhU/pTbg16ni3
mb/+kcjKBE/qXR7SMwJ/0G2jVXQz8kMX8sC0Wuz3dqumHC9TbhqXqqoSIZwS7mCTLJKdKZ/9VtJj
p4Frgn1tTQeG9hXyojErm9TC0QNXukHRTkLjqFjh8G9OTYM/hnCH0ULEqnbkKY/vZAqd1nwqPpp7
eFEYhbwaDW6TYje8NjoQTPkoTmvblvShj71wgiKoGEGnUd/gmHrIYkVrM97Qbikw/PsljbUZ8Vpl
rf9ONyFGJuLpqkdJ+lKIh5UwXarVYx3itxexK/zR28aN42itatdWQw/SUWPVwwPIYUmHmsS6VnVL
panmjb+fseG05jzcajh9PcIZF7DaYxXMqtVRkZAO3catlAfQ8LBHEcC0MvbePwH5V269OTwbl2dP
fk+GbIMjazLmtGwztc+19M5jCYKkljF3rha8QqM8utgTP1zgABaMmYkq3DtL/iCpb7GkJAw6UnUO
XQtoDwqYLuZhH+PstMKynQ8caFT22vV0fvqSqWDs40PqXf+vOUEoZShERB3Qiv5sbpOApaJqG4/C
3CTDUsnr0FNJVthRMlDmoDwi4BvvR1elfETCQpyk41HEbf75ABya2gYaoufRNyArrIhSbI4r+kc3
nq9Mg8oB3M7UKHRATpU3jpMdIR+EkJcj1aU0a1AkOIAJnqXN9sVMHkW5rMCKViQ4wd3W50wlWtjM
q7722nn0UMQt03MwzZDlo5qlgaMW+51P8PRgrfika883Scq0fky2rqrNfsbe5b1d7+Rm8MDMrl1b
pioX0mNSJ4HFWbEL+icJv7LqCIY6L86sbj0cJ1hhDB3Q7/yfh5QSkRMKQPR3ciBvLCa+Zye7HdXm
rivPjGsmAnm/pq8OqJX2JTIJ8Dyj6aePetTDz2Um4w2CggIwJnHM5fFYCvkIi3rg4lO/rpqreY0h
OLIFMzHPrPFJI+42M3steLb5iW8EVSWE0siqEMjXxw5vzuqYKHpPe/YcIXI3lVENWhpQ5AhrfaqV
fkFJE16j8kxN0ILcrKGkp7AcP4InM43jWv9UR2k2dD+2vqGl2BFBkogSFgwQukFfrJeyCpaQekDC
uOziLjgQvKqh2Ivp7ChSwc5vavSuYa1rfk+ovfflEhc1r5JmfX1MrxOuVrl23vBoyomvkA8WQx47
cLUjuXB+vYQ/WfKI9v+c0qI59UcQzFO1K1giwpE32pSDJDNQsRj5GffI3g45jby/OUdu1jzkHCr6
fgJv4YIXeW2xMqzCgpjSTbzC87w+LtC50wdO0NoVdmDgsGFIIYH6Mj0AGWKsXsXI2z8oS4BM65s+
jvbMMhCb2w04xsPRik67G88Nke6H2dlTIXXrSgu8vA048aQScb7S94pBgzWUn2gFNRmD05UeYjfV
ykCCrAuZdrPXURv/HktFBOfNDGeQvE092xILT6TyIdisPH+ImczyY2ndqVgzT6urxVK8NPiHjMmT
AoXbhr2TRvdPKfjQxrbci66L8DDDh8H/RZYQ8tCuGFf3QGDll0xbPEhLB6rb5ExRXzFfMfzGnARP
O91hTOTsINXr0gk6PfLlcFZIMRFG+McwrvyiSfgGeNaoQ8/+ioXQAmIvbiAr1eq4ndcVNo1vY8+O
uwJZON17L/kQE4xQyMhS1C7shnydiiiK2w7nBfPqHrr23fzNXfT9g0zslPM/QKyRN90Ny8AfJaDo
ZJxFhzi1dLYsYXaLFjSCJcgw9e+1DLDz1kWbKq6CDUf3nl5MF0nOwi02A+9ces78remESe+4D69t
Fj25AzAXQ7x6oh6OYOj/G0hVeC+Q1ADegutBvFDAumLEMFHTXnI3ZUG+Hjdwezn9OykeEhw9lUxZ
lTuoHr0FVxcaQVrPX03gA7dCtQIhldreRtVycu9uA70qEjbGOEaf6Nus+FA3DzeTUsZiz0/UJUrj
45CrRSyU+FhBcaMilB0e+L26+plcuyoCz6m/vBOip8vyaD+ku1afLAyWfzipd+sV4bzaNRs38PEt
rOBlWHWUqvyhXUx7TtclKvb0YRiPeeC60vlT7dni/9zCqcv6SXOTNXoPNPV2vIyZcH4U0eDvsWEN
/AQfvBGWBJVuSbZeEZ8/0aAL+xRMtYPaAadQdUeuBseLtZBRG+qUH4U0R5Quxfw9nOHUq/7xqDru
LSOI9TxxdsBLAhONjY2GVZaRFzs4NC5iQsOa3ftO+jV7CZfiounlP0bgGME/X5M8hIkQHP2H0LZ+
HhVSklaPkCZCs8bYEDw+8p53vDf81yNwx5wpTKodsuJ0bvlVBlBJEMUbJgKk8ISAsKyML8g3gK8O
WjTNYo3Scgxxm8k4drz8t1pO77z8+bWKOIfzVEqR7ttxpd2RQZjFU83hkb6CskDTQgXc5jJZ6Kgy
yGJge9muytMQbydFc7wJTRs1b75o3RMyvJrCoHrfJ8Vd7o0H2qxRB6jnBd6SNE7AAx/dRCskwSEr
LfmCT0ZUp3xlIYLXjN+xD2nPOGYp68t3XxVcNbE9ucB0MpiyglWYSdRTqlcynEt6Cm8/pciwgrXG
lRmNg8F9AazTfzPxArra2cRMPdkxuBrjYOoMYsWZOq33GADJV4CQHTwQHD8Jg5c5aI/0Xn9fAU7u
VABnzSJMWO2zg2iyWTnJYLaikrXpRtNhkAyMiZ0wgSV7ebsgnLibkb2g/ZJds6pp1m58Gj3Qsb6W
VkSlfgxUlY5kVJd1aCMMGKY0pdvMM273o3pI9zOgVwzGk5/SKvcmE11lCQmo3DKgMYOoYny8/tXR
G3RydgZ4f2IxqNSif7FkflM5eOGnRP322IsrN1mGTJLq6AAmeEh2Els6DilDSYrBC9fdT16wPXoZ
k11dzBU+Ym0nY+tkjS2TA/X8nvhvSfIEpDEcqhYN9JB4BBn7uf1lYakp8pDMm+Bhu5+TvoHBHTCh
/9K31tPP1+MvGvujhFAwNfAXNHC5O7xVezVhSZcxDGbSpgotZxdB+6o3mE/w/59higQj3kjhHZip
TJlcP2m/hIXZxoO+9HLBhWeshOSmZsDU3YaTOX/PtXgmirOahuydCehSvYU9Bm59Xk2xQmmVcRLD
DJS4ycOQUJ+icudyuOyrqeHOfuffNZNOFeKcENk8tSmzXK87Jw4LKvSVR5GLJvwvN8McEKpselV4
iKXz1Y9Wy0dxaL3REcEwZbdgA5Ago0GKw8qWSNVqk4Z8m+duOQ7DwWG5JiOMJS4AbXDSUHrU4Jj2
/NfRs75X8IugmFcNpH9jfl40sZjU5U+vXCGhkQ+EytB8+8FkY+8isfCbv2UaUeHx4WKvCDz3wLh3
/o0IoT4On66a4E7Cg5AUNW5iP/RUkacmEnJeg5bDL5IbNQKa60X5lCkPTojWoX5mUx/2onpD54jp
qh/m/6pTB2mmpRbZhyZiHx11He0rH4xiqCOwlN3GTiQtlMdiklEsraafv31Prmy/tTb59MMvlRsa
3n2+qBuRLLwlccOBv5KA0Mmsik6RoJ2cuHfoCfy9lwqnvyUFO9wTcjScVje6s4VRiht64ikS7Olt
U57mCpiHD2EsIS/LHMCxNjNr2pshYDsoaLVXwLnnuORo7NF9+A+XN2vZU5HQcTLy541LInnaCNu8
VRhRZbTJfMKhi42S+B2148MmRtHKKfCsr6WBdjCWNk2nyC9Bg+9Rn6/Gz1700j+Baf3l7nJhZsA9
BJCfV/odcEavh6kkzPhCGkA7uJQwJVKFSU6ncq8EjDhEO5q8evlf424qF/sKbapMH3YJ/4YaReDq
xt5SGGFX2oHL76fETvs7MKdz02k4WmoWVlUmG3ED2QgfDWNEDzBDiGplAqXz90Jud2RmVSQ18iWM
rY9vHL1IFBPIEqIyojVS1NMUrpHbCVdGCENnL50cT4jbi3IAyDbsXy286pcZXIpIeMwAY/iTrvbL
4W563Ffk4tfcwDkhkFQ4v21uK3+3ev2h78+OAN5yxwASXQ49agjOfkL/nh+OcECj7VsEYzdXWKwa
OLT6WhYwNXswjeYTQs2Kf/cSZtrjYaoMhVOL02RVj5Xx10IUJgU37VTL6eyVgnI8g4Pb4ViXqIdz
SAb7Q9Vw2ImVD2SP2yxzxH0Dxe2jnPe2TjIRI26pAdScvolGoyGhZQNfibJjUd5woxonA78QDUe/
XlCDFe6XYsrE67MOpeF+TNzUV1ZuFf+5zraxkpqggwrTLyzas1C+dtal4qmfuINj1gjAp3UG6e0m
F3akUonAKCmzq9awSTOBKQKoYZdtfuIl2ZYYAsSUB38H3cLeMctbucJ1TTdytU1y7H5fC3/7M/IS
SrKckYbMtaUEAI3+QWLgGBsCwM9F2CP+DJkGdNK6NMsTbM7Ib+I+AO88Q3XRiBwEGphAwFperYPP
/7ptVAEX8KMJkFPmovA=
`protect end_protected
