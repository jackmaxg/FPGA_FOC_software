`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
KrejDm4oONuYm6eoIc/oaYTMSg2eNjeKBqda0EjXHPkR+VoMF4PriNhaDnsXF+DyTMZm75V+RuD7
nWpqddQ3Aw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
L0sPDxM09ajABQg3R7D2WQO6pfG6lvfTeBI1OOkv2/KEHi2yB5zNP0SkPML2mr0TfN7jtKbuk5Jh
4z8voSkmrHitIaXM0NttJNAMxNyKUESr7nyvNGIbv6L5Rg1xms7jSznlVehCqsXIdT373eQflR+9
RiY0VXKC9SQASFbhYc0=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nwPd/kSs+pKxzqbzKrG84aj6Lhs3/i5NLOCCpYrLPG78hVmy2L2n+nDg1AagmyDAd/XzNX/W9lEK
rRm4FL+5hzdV13dgVeMFq+vM0WZmNBM5+a412h0o16xdAJz11N8zXCnHIU/7fDWz7RJcl8+owt9b
yRbbsnH1kimhNdFw9dlEKCa5PhK8Y9NjpMQNhsIFDugSHtxlT/f8b7xYFp0yYtoecjR8U4c6DCk5
pHB/FXUAYKQpbwbaSjU6hLiX5PECqH8BFL5CE5swQgIq4EHgHMi1kpvNm3w6IZYkK1FPXUqne/Sp
z8KN9vIWGD0hZTZ5XZvegTQuLnQGqRCw0CdnCA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ByVE0Zp6xXlrjfjxHVTbU2+PqPt8rvJ1VMPnKfzfqMYdBDpgXAKTdNQRGarKJSOwuEqBPyPOiGi1
K1O9VuIy2Nn3rs6rrGTfI/K0vasx1+wuXYBA2Rb0K4IWGF4Fr0C+Wt4fRR1ZrH4XcQsEyXbjz2tU
HykeXUzzU5HXxXsbSTu3My0gQFff31qo+jul1mwIQxGu5kk//bHHYA33P4hmhfvsQq54d0O8HzVs
hoYK7psbu1cPMMyLTHSw35eFsmTpYMnZcQkd/WDghuEaX8KQKYWaR8E5xSrI0gRO9wPLZMNA65BT
Es+yRhFspdz8u2T4oVJ1cx7nWG7DgCx+uMHO7Q==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
U1mdpeWGlSnD2kIq0uZoIf0/FF13I/8zQSstV1pkREDUsUsWTOD+VPBvAiUg+bqu4bKdQUJoll5Y
L5WRWCHy1GOhrhcTV3NHbG+aCmHA0DVrS5+955Sp0TnUYzUyWXy9e7Za7eo4ve5AAST2rzkQlTQu
Axgz/naoqIcmpcRqyrN2uEe2qzcSj/qeC5J51VvKQJKTIweTR8SzpHrT9csD/j13Gy2L2/iiBwyM
WRmlePefvLLiCCAcj9eFe3EJ0O2oOiKoUdEdC6+96sepmfXdDEtJ7z+cJVFPwwAlKpUcwB4xH9tV
lrcgPPgvGarP5lGTDKjk/NEiBS8JUMwdNRfu3w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
R4SJuEDUHh3ETJgxZQZCtvf8fPjYXlzMpLlwfseEchFX50gJXo1st8+d84CFiK1N++VX0Q8m/AMV
06jBgNJJrpWqNLKXetqTdCLakIwRckeHlaSR4tifY+MnS6hviYMhnh4s2cueWH23zpRNN535DF+u
hi+wuwR5xR/rIZY8ZR8=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MSS/YW4GcS4lNnbZAeEO7AUPTrdvy7pQ7mhHTgW2y4NLSu7GT2Er0v2fvmezqL00SfEoUnKtvwzO
kLd1FVxyTiwQch3y7+Mg39Wez1xgLz/KzizmX+19T3Ptgs5vX4h/CdaxNtsbHBvhO78cVw4xiYJ8
p70tNk4MpfZRjPCcakKl/nvLJZfeGb+LZIr8i3k7TxC9/vYfAe6BfYZipqtjgoGeQ+6643JY3mv5
Gi2zcceixpzOaQ25L/EojJN8CNQeTa7iykOMhnZfVfUGiDAu3rwyRY6Id/+qHIQkOD38e6xEmrtm
viVcniQ61f7+uGQchrKrFf0FAwdSlLcj+1KW+g==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
phEOp+sc8X9th3VzDtg7VdM/UOq2+wJ7AfBanvGUq7mcbdr1su7Aumludr7lKQxD61/T2DzvBePm
jd45mDc6r+LOARyhTuwJ56eWr3jgMqTr29XVqMkKntPJuoF1nAAMxFBQuVo7eYFoGCNya++nkpoI
SRfCU1vaA7QVJ6gOZ7OxJnT9D9+t3We/KPufxAOu72+FetXL8nnLIG4nw8rdZF755qrj8UeMZiA9
rch6twJ3VgTXOOz9cFxgdcGZHtVlzvwYwiSTSRL6rh856wioll0XlkqAoR6WBLbwTmkvkd9Uca6R
pC/V7FZvZHTXIAVR488nvm3RgDpnGaxEu2/MPg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 432800)
`protect data_block
O3XXDYbSEab0ZJRyaWVhghhxPmoao2UZKwYNb/lJm3folNnmEdgTUtu9e7Uz9CXfToGajCTig/sD
juG9W+b7xyh55MgfE15obGRiuSikES6RivXWCZW9PYgS02MolqV+erxR1XyPheHkn/qgSP4tzEPm
/e06GyY/rUWLmPJQ3cqH4HHVXa268BYdXOlBjbVtYpXno5r5N8qFls1KznCxZ7G0xVLb67Cyv28e
JZO9hyL19OVC8+enRrrjCpH+ERD4DDrEHLpUH3AoJPw/M4LKPDeWN3Tf8WiKxIuwG0204DXE8S/F
wZJt/M70SPeWmgbEArS/B4u7/7RT4IEokX/x5TT9Hdbol/j5uXdCLt+fpIAhg/8Ol6dcNA+fxoCZ
K2nJIUDlEdsWWELT/nWzObALQb2iVBofEOfweUIem+HKs/7W1Z7eIIDQi7Ymv0gRLdPG5GN3Owj+
TteyA7JpSepCfFDmIp7Filjgq3S6PNeQwxQmjuloieraH5KdO4yWnokgmT5KOnoo80qDEh/zNb+O
Yc9d/3gQcnYMfDn8t1+XPZJh2dtz4rz8ID3IZWkuH7OkRLSo3DYouY8uEFPdXWFJHsepKzmQwdkT
GR8NpL6O1A4nByA4xnlYxGZhgnEVYEtbSMJoBmw52ivSeth/5nad4jxNtQFfzG0dQEmJcauQb39x
p8NCFikwVOUUDksvQHMpCZhDFGgzV1Pf0vxW1MXBAcm3uLy88EZxZ2EBdRvq3cyj8fS4CpIjUWdl
uVcJ8Baa8FLYBWUcS3YD701MYHO/BsS4QxiH51LhbfzwjhiuBgux54A5kHiA0IMij8i8c8Fqfewd
NtRQ6iVeZihGsbYKLiaP06nCUiCenpfmj0EwJgP6uXzQdbVt4EPDwYKJESJi+vsV72jQx7CNKOwM
ZHYj8lk59FCydYPW3j/UhQWF+7xiwnnalVJHIVNgHK1F1Bvduhvi3SM8hSZxpc4r4e3v8aqJKYNg
aoYwTLywSX95ok9fU7S0FmdmIb5rphM1d+xCM0lghr0n/7B8Bl+QcxB15NrhcFD4c5twZiPWE59j
SXvaskrjxBrujK2XytpFC7XSDhmiMuqCD3ifTEcKd4DDCCGypSwwG1liRZlD2ACSXqSPRsZFiUkW
i8ZazG9yZwKtgbgrK+yOQt9gTcKo20aOQ+V55rZ8uAt2NlUWKDgANfbDTZdrA2+3pqIRqEQM0J5f
5u7AVe79xMiQyiioDaPMvmX4OYS0GmwC00Kip+hcVwPO9Qqp1PyiK7MP0yMqgnYNEaZ/NO9Pvy/Y
r1x3WO0gMFtXLP7Tz7Zggd1ycgBfBW/t2GC3o60U75atxLaNGfYz6U9F5As9HxFZgymTLN+dSRdm
7eBNfG+dj1mcFW3httFyNhIaIWiXbLzlTT5klggpwgpZKBr4I6h7Rl5ndxD3ihP8OZ+6m1yfDLRD
toahpLjnecIbSceIIDVBqhvQjvCStHIQ8RIWFDIsHMqpNWWXqJiHvaPFKRpc9Ewx4beILnKlw7x0
C+M2Wti+++j3DmLMuRLbNrDSIOfK/DRWBw6+Tt3A5UIAXyQDgZ3Y09C1+ulh9gC+KSlsa9Yu3FFX
E7S1yIt8OpbFUs+ZMyrp+L3iGL+DEbOyP4FlkwI+vzdl8DnuiHTZY7zCUYToRjRVCfXUuonb1oxm
mTgy+RncjRQi1o8Fx1cibPJIDsksQOzwDpVGvBEMtxhYuNOQ1bXq0wAniGC+i9b2hlt7RCwt2jpE
nqKN+AXjieIzU5JaPRMdEXIP1YBc1YOaphwRDFxJs7wrhL+3EAqB2DiCNpCjEvBiPkjPiO2sa3j6
T8zAxh5NlBlUWohGal/ucLeZDSYS5NLmmQHTvxcWuNwJavKCfRQmr4hnEIdyMoor/3Wyc1Y9f1HS
O/zJ3ofbiKli1ITY/DpDxOLgeLTZUbsofO7w0rDWlUeSP/9NXMPc8TvwnPtFD6GPQ/FKdFegp73E
VA3uYmmNUSUPYiblhRvime6EGRClam02plm7q+QJQ1dqaCLtqP3S4czYLV35LTNS9PIwuvh0B+di
Ip0+6cwLob494ecH3+DsxcxPtkfPzHgEy9A60iCHt4L1t0WJh8tQbCRxmgWTVLflrc/+LndGWaw/
xGKvaLfveoeM7k/zaLJsvUzp2cfCmL+AaMii3fD5sXPgzDg9eLtB3EYknNaDVEQK/hPzqsOeZMfH
mgyuhM9UVmQQNvy6VsdlR05bZxLWNMAKuiuStTzeIwzuFgAHyWEcf+9jE+QluXADOd7tyhl2ftJR
R9PZ0b55ZwNBr6ZvuNpsMMS3kQZys4BVPTNaEzmWJBjBxQ77iC37OIN7h9FfH6kPRnhHkF++GIUU
0sOwtoc+KTZ+hWsOKi/F+RpiW1Uq/ufzdxWu0rKLio/2afUZrwWdHLCST/ik4eW3zXlZkaATmLZy
P9VWvfHIRqGI1Xh3wwwjKH1xoIqk7SNZH5nvQS4SGErfbUmH4E1DOUH//H1dU0LRKZGRbjTKW8E+
m12AqNGYwVt3Yty/2KmUCvSz5avYkvuBrfY/g4KbuoIllX0ubybsj6WTIWDLaEumbjN6gTep8kGP
VMjcipjhy7NokyFDEFc/0kcHJNb5cn7zbZ5yIAfBFzBEkZzpMIDXC5ML0iCkjzT29gOy2GoY7cdB
8N+WkLXeBgV32oLzyL0B2A4Jv8u69jJk4+xNhrm4uMU4O6yZ0Z5ExFGZCpi0YtxXt1JAbhwpF/hF
hp5q+PK+zzH9P4h6RQLHEh53RHVlVXPuh3vyGR8RBy9tXBIIfdma9fM9Kqc5uXwefFSGQGJXallk
rbXTGwDBW6nB/TjbpciqkGlQAat3nCyc1tfHuB0yP1MfOTy3cvkfHWnLv4k4U3OeDtNb1iuUWuGh
Sns+uXxiYf5wXArBBJ/mP/2lfcKIqRvM8B65iFSKp8Q7gxH/aXlTqHx2lgMfBYSyMjIHuWRtB1up
DA/bgjTTI/2e8uVa9mRBzjDPfV5ZA4AVtt+OoASl9Y6mx36V2+jz5cYJBUW5olnAB/agmPulIS5x
4XpFDBTTC+hMLZG6nueSGtjjuJBX0bC+8vfeYe6P646691rxB24O8d7Bk7qhLSTrRbrZtq6AzQC7
eD+O39WDLoKY/oPcdgMsosctavHkPoqHGsBdvCYNyN4/fL86+ozhctm9sjy6oGqin3W1H/KpcKrf
kkzncaXK2CKugmM/bep3HQso+sZgHMxXqb7p0x1fKhDNTH0XSdcsU4nQQW2kfNV2vB4Jytld8+lT
QLOW5hYV5OHQcsX/vTLkxnkAAnDETDOtl4HkHokH+vNVVWXVoeUBwE0/QLuZ16moVfwCBU/dNkdV
i4nxMqQrxwTNYuEI5Mcv0DWYntgMiUSBzfIi+mG2D3OCnGkcG7DLvP4FIeGe7yToi1jBxiwdhxF3
xLDGAAgUo3BsgqgNuespXGRvF78MoeLq/A2ZqPZlAHnWLvrV4qPfwb0U/glpnsJe9deMfPW2wfH3
6/EmPk4j7dfTY/4x7YI8dMaX8b89bo4iOMEtXxKS6jfl5FNVREwPKfLp9U4e8gWwBmOVqMymYQka
qUHVTMIUS4AvlRoOEcRi6LemljX0sEiRR/iBoPAxylEyI9mYzjYRJlLy5IyV3wCAiBomxGDHF7Ll
HVNS0U9NC9aWR39qEoK7R5Tvj5ok93g87c9zYk31jQe5ruAjQDmqKOvO5Oc18RjaoTs9tnZ6Gq4F
3f3ydkXy9fLNbLb8unusuvVhXxvG2oQRkoa7ZfQnj5tWCjoKhi1Vrweertq8HUSOArSYS35JefTs
z5u932+TzHoqIQ8MyFtYC2+rrzLwCxU/7M+rPtRDUKcIWG1vXsQATjAjjQCSxPZtmdbt/ijnWj3H
mo8aaSxoagmMBKfeD/VGCF03XUE1hx1UfYFP4BMnK4IU40iL5QStY2bKwDFonn0Yk3sy/2e8V3st
5BFmL3eJNvLvh6noV35xNwoW8UzMfNEWe1M5BqCFYFHwebhr7xJAtL6PnOmL1USaNwWlFNx5PZ/v
c2w3cWrRNTAofpOKVZ8gSel4UlWrIc5KUKw5NI3EaKByyLvssMeEyQu5roO8iv/ae6wP8kLqBB7Y
1HJ+AYUDw9g7nhpQenvmPqaIq1CNjSvVZtMig3bBiDh1uaDWbNj41lan3FEbEkK7z8ajXXysULLV
o2/3XmQfWdF0svBqR1WwijO9lcqUpa09ToPd/nQpf7lbblvndkjiTo/GATmWiDQ8vyUWnOqBo3xP
zlGDVXw1c/t7zNHX0d0H9jHDvIJHYW+wiWnbYNdCSTsUnx8Gxyz2Zl2C1vHwdFZKBD9WAxdpY7GK
J6k6zAutZzjxI05Z3jFz+ogDqp2huh6ijKtm0aZr47kk9rNIJ/RhxO6kS/hOzb6oawRgD10zhqJz
qOojXL734bjfnZcglTzlB6qMW93BbaZsERSHs3Y+6SAfyiBLx4ihRlwg0P1xV17/AwWwm0FGW28q
OcWa/PIgGsh6ATAFCpgkBHpBCMwEYvLYZNqPFHrOptD5xWYOF0hq6Jd1sblBGPejQFr01iTnyNKU
EhFEOHCFO08lPc7/fxUD/NqLxQlN0/MfIqF3O9jnRk74iUzKtrom/lzdAhKmvz0jsjmONeqUwt4L
dLBdPnwM0H/K/0jnKqcbXQ6M3kv+eXFVGiNIiSdMJsFUm8ggAb+vDoPvWdmV5gR7XfDOErwXhxS6
mrvoHAgjc5Rerli/Wm8DojJv74L6lmrDyHb1467xFrFTJymHwU9jJVoXMudW/CkvOD0QHuxBOekB
6wngMYPVyWWu/CTjNIKsB2Il5LBueDENtsLF6wVTRviF/mZxHsq0eTfify6aWAmsLSGOkriiyGx6
iJPLDKQbLUgUjQOoRI+DsnVKlelzjF5mHAkoAICQ5+19wshXJLAy0VomOuRO2g/mo5kHK1yCfqQJ
ioXzdmWqRe59agBO1lrV8p1dfgmepDE518WR26C+PICAp07ZRpJvtmu1tn5vYbJeFJ0lNRVXPgkM
+MndkjxxowALBgolUHuQhs2gG/lEjHiATubh0zt9JzmAZV1raio2iSG58vj9ZCy0VPEa6cYQcrMC
vWRlmM4HWMVuk70b4cffBYE/I2ngd2e7DV3sM5v5DqFX78uh65kbrchjFpO9S7aIo2bLe0QoS426
tM3rTfrw6e//p0NEXhYea2XtbOhCSo2CnwTyHovLsX/f/jCFWHUokzyagr9gC2xZlVS1z0Ztt4il
YrFkLKoPwtvmj49uSmFA4s620hospqLRidmwcqzzsQcQQviBbD8eIO67eZnw3YE/YMtIDfKL5wBP
COJG1hVA/CBl0mgZc+0IZghBObUMPs6nUjihMSwVEax1p1+IUqT4UTEWqJbPZZ+9/UuCci59SldJ
W/2JtDDEZEFhXiRErW4THHGp0IoIsy5qkzoxLVME4uQH9ODqbkhbQ11NLbrRwoKZ4lpCazMHqu4l
44ol/o4YSmR2Gx2X8jAW7Lfv/NZBl+hsgKF1f1Q9rfm64L9ihUXIFrQchZd1bmXe0X90ouI1MRDW
6XWw+y2ZMM0IGSAnR4reAuwBBmH2/2UEV6cp1pTfWE2/v3gwOuzGkFTJL6q+AkQ5Hofvm+O3Wpyf
BzvGdDByJqVq4Rpv234+uOGIEpq7Eno/PLO2DzIM6CT+fxgDN0GGx2md98oFfW1oxN8XbCpqfHgJ
Yu3itVqQ7+x5FLUXzg5voO+oGheaNJv+npYsDgo0cuez8vNPhaAMlerEd15BB3UsaChpQMohVltw
2kNFFr5bBtYU7n3HvBuZd4c1gAT1MjBge8I8y+9r7c9T1VU77uQ2Sh8EWyOzN+wNbbiYWH58Mltx
ltP9jyis65PXv6XMVX23OEOdb9HcAYBU4CDQFzInjRrsW11+sOXa6RNBfOblx/VmHrgC+jiW2sTO
dXFgVJ7xsuNtM4eO26o+xxeWL9dD0Ass5UZUetBBF4UGz5Y9upTcPWhtg6usS8huoGgYq2sMwBDn
8cVWpPprKpNLR8UyWmiB1gntflfTjHXPGiR4BxLFco0QBWIe7I874eWSAqBl1E1oSQDadLU0R4Xq
Q5XGRT15U8Az1WWvt9llIW3mfHQcd/mgcNUlYTLxozUi7XqW5iGky1/UNDS2BUhUOdh0YKjmE+jd
0r45Q5MoHjbrb3fW6vyAtDC1uRfAP4q7XF7SNPNf+5J8dAih15s1xp8hX6dXdRgGtT1hPAONHufb
JV3l+qHW15e7wF2mrySEWm1emGhWw3LYEXmmNANsnc7Xi/+XxAgki4CbDKtDfvrZqR/PiHnPUI2A
xE1AWS/U8eCxPZJokehlipx225lLe4YrrhTFZYK++MNNOwmO2PAkzFFnYYwQ9ch697hviEr/bif9
ly5QUuz50Bf23hlLk+ecCFfGKOMuMpPg/nftd0K7qx8iwyzXbO+HDecpyxvH9MrKjmVXVAFC0lCB
Cp+Syn1EEfMKG6goUnWNgF/XPvAEdqENUaxI3cnxqG/iY7W+WYhqWnjUFTlA7J4BfeOfVnOmUT3q
fVIVAiGrYZNxwuXXBlp0cO02L5muoE3bop/A2EHuX0ZmUvXmAYSSXQjmxxkq1TQl3cGwtOpbKIme
9li7Ck/YvEaZ1hggHjATYTLVzvj7QMXfSEBieCe4bIKQIfcrIYxyrcZlqk80yrXx0bZykjoS/Lgh
Rl0CjNsvEZ/82WdHILFbrCnh/VnuJPzrPsFHjbi3mfW5YfGqby2zFzgw91piH0ssafH10YJzIA0E
fJu9SwB99Rg0sXyTno0rIhmA2n/jRRrF3IJT05U5WiMyX+mpxAJF6S+WNU6Ic+bbmpFWmDM2yiBf
NasPmLH+8P83Pp4QAcUPfJdB+wPTuNuYRgIhRmuR+bIzm1OzFMWatXpG/HKzezHUjgDmDIPqlmPo
n2H0/P+6lT8M9uIQyvCW7nBK05vMVYDG8deNZCIJvmDpv2LmulXVq7Mg/koEUYEQHrU05TJl1vHV
inDtBiaJ+IoTVfnLZwI89htA0kidbyHnxeGgWzEdQTwcRza6EiUx3/JNZjbZu6cMZUPjVH+ZfPD1
M8yQxjxxa2ywSl0R2fJ5P5KZ2g4SMy2YNQen4oBXa4fvYFT+3s9xbZjSbJFfizNRlsbqNzKmOTi6
YZOtsx0OYTFWGc8WeGWIlLAU8Eiv6N7yEVX8uhO7qT6oJc3AYiWHh5MtNThnx+8uTL/C5w5NFG/K
Q5V1gaM5l3+4meWQgaigSBbNU/fSNmFZ69eEDAlp2KNPW0uWhwEw/TUyrBX6f/oT3IcLzpTZ12xi
DysvsoYS9+IcxSECJgzy2n6NC/uYXVg6zqqLpnNPZySeKeNsHIYotpmJH3YJX3JSe1DUNYhf9+Ae
O1veISFLSEzn3VeAxiHr/sOTrLkhOCgjJ6qLPRWqsdEGJWks/fLmZuhp2S8qPO2FKYg9Ld9vRq7K
Zvn7EKaGAGYpLXAKJ4RkRI1aH3MLehAJ+G3Vg5iNL4QDKHaiDEunAc/1XU349g3DWfcGFziIGHYr
f4nCIe3DOvGs7N/2CUuKERmL9FFh679cMVah7bkZD3z9UW8OQ1BYZsiMpYwroHjse7Vl2PjiZ9W1
b/BJE/tr2nLTA8DzF5NTZqmgKF9o9I4FnEIDZLZliUSA+W2HBn44OBxokbj6V7Wt42IO8w6CWboT
+R6S0D72DcFeQ5XuaEJCNSYs0/gczZgJk41pejyF/MXtuoT7FmdC9I/WxK1/UMUNcK8TiaGoGiGZ
rbJBeQtk57wmeWbxvIJq/+cX2rX8EfTwhtAnbSMNtKuG8LyyDsx5Fu0oVWcI+PnLUzoaat0LsogA
6uPk7fNK6wdBhQM2O8mNeMnGQ8JdJWxArZgaloy612wkAM3x/XllQUDrgZfG7zIR6p/EOtFWfwxP
UHwAvyONXbtFEVTzEYbrKd3mDJybiYrw+ROPZG4qMGvtyMKFz8GY/h6SrDY5DFIuTOUCMHhhjxnC
4txxL06/m/hWV8pdJwhM5ncAnTZBBYYvzZ4IGPVg7FIkei4c2Y4gwiKgHICSUVBqNxS1k97NJ0Mc
kpRAiBwe7CZvuEyaP+ifcwfyYD/r+66uhPOSs/ssZU/bjUp5tl9j7/e0mm8+oTEh58HNkYUSauri
V93i89TYyUolrROU/ijcbeP0yqOX6jXfGQELu+gwyIa0bjcD5gS/zuJgXj3z9LWxQzRnPKhs0Mtp
T6d9VcyQIh87tS3y08MHWhaDn2CFnkCYtdGs3zLXUM3OCFP2wkxQSNzgDwA24MXatPL96i5NCG6u
kPURtjPJ+f3RU81OU+1usPg/ZTYh4iAbLLPEHQHAC2+Na9EhynnHuLPDa8IXHh0l+MZaxNP0hYgX
zz3XxzXx++uDgVZl3vUK6EFdSJ+MJDbSX7Lfq/tHa2fOCtbdc7FOhTb6mUfJemLs8rVWfUklxNeU
2Ldsfyl9zMPVfaZLmOZmkTghW81rNDXl2HBGjDlZRsIdc8X3iAthutjDggTym+NitXSfnZlwmwEo
ttL1s4AVZ8UsBq1XsMlECm3IjqJvXTu3feyo/BbF8/SJsUIwDRtrwTzKgXlbMSf3HZXr0obY0mRU
RBDzLSMwA1VyP6c9zsIdG2Hf+9s1DLM9u0SmLGsuOThWqpZWNxAmcNAcn6KMi5ssxjR+omMo1geH
HOvFDIfttLVQFR5dW9C+W5l/f9l+0KAU07yKeZF10TpTuw15GvLpAxRVkmuMvPpj2eyZJOBMxFWp
Qrl0PMrKLTS/JjUPrOVoFvbM/CqFArQvkdpe8+ctUORM2c0RP88SBNscxev++YrOBZScmqtdCq8y
jcT1p7sLXqspD5fTtMGAJ8vwxl24/TlDtwiQKz6OawgZ0gPX9MUVQDrU3IlPJkj1iMTZn9Y4O0iu
FelYRUjRsAiSnoOBmD72jmvgr0qAXAYqqWwyOxoCwDXIGhIZbX5EFYdOTRFDmAEQjbJN33fUvFeq
WpKPIwUrZmUw7gZ4k9Lk63DYDKe6pSQFo4g5vwVCaWIeR7pHVDclYW31LVdvchaAzGdD183T1jxl
n6tQcIj1SPh5hHiJPpnfu1SYh6hGy1bcztOvEDDpZJ8y59t3dmtdpNe+I3/00fK3Jbsy8cpNNGVk
U96DXvpxYTfn5J9JOf1r6DaCy7Ztfrftzx6uxnSEvmakcIG4L5Q22bnQexL+0NQ3WcMqeBwMNE69
R78Vvb6dLs3E0bJp7IJUER7uNMjcXmkeMltsMt4oPOKa+KK7cZGm9giX/D4LZVH7iZyBniRF75YB
lMvK266v1dPu4lhOdpkdlgwSczBa/EJnPE9WEpWJWjxRMFe+uajQ6ARyCJHCPeCV6Cabhln91+XT
02+PlTGd4qOcWvfA0fg51zKzHwH1TRsL+2y3DYWOY+BGoqwYJKxRffzUjSx1z/q5S4BMijfVTYe6
dKyaKd+FYSBgyQU6DvMUftgb+UatuVaoSmqLnRADLvWsKFFRA6Dk1ENCuhettTQPD1hiu7/Bjlr/
IsF5xlBDTax5zVB39gdccfC+6Llekttx97pYrs8RU0kma2jExX1gyko6FhgWmWoRI8GBxthm0LDX
+lI8Y6/0pUx4aqK8meOlUn0z1pRNvWRJ5CL6E545rVWadIHKRuRis6H3KOdKIw0FIVNql2l+aeHP
WSN1u7NT8rwZptr0QodRs7ew1BDk/gvB1M4g0ypG5cRXMbOfkB/tv+BuNwMrdlAq+9n9MWYmX4vH
wUDWpqdpM+1GCvpmUfVnnbOXoJ7jmn0VyX+zVehFzgBEG5oK9WtX9d3jYUfQtyiko/j1W4ttM+fc
4sT4b5zzM7B3JqDyl1N5cqZCLJmsSmlSEbiwldUI1uAnfxgpWDSEm2v5Jj0mA+3lmPhPdaAxjpfL
x3I6/+nmZw7+Bk0QnFVlshEI5/98D1xATGqsAE4Gb3XyjIPY8tOO0xI5MFiywHzFqKzfwmv6hwcY
/m9R+qsg0JY40lnuOLFNCAgZ8aPrIRdUPSJjC7DeaWKttELIK7uFOrRofLbRu0LGkWEg3rQKYWSW
/c6Tdy66hbaqQzU0BU21JCSVr8hElgX7eisi/w7EVBtp3roXeJinzbuulKK20LL5SznruWaa2XHG
CQYllr8XIlaAKmt2sdZYl/NnZlgykTzeA1boPTQh7BjDCJD6/NA9oc8Fg34JUm0II5rQ1n64U01q
5MBusC8mV5LwaHAK8xDPB1MIHiYsVpF4bbninKt179g02TN42KKlKy/NXtjeG8qNBhBhKQWzlsPT
J/ldTWyy9ZMJNqV2BfBPRXJcFHmesEd+Qj/bA4Edwy+JUNdhwV4ThevitbzUWkdhOBiXmZxQKyL/
0JDFUBlhrIUeDi61K4Z2Ct81g/cZOc4yHrZiYkyWQzYb1IqeeHE2bd+Yc56J4g4XsFtqKBfFLirh
Pw5Gij05Rd0x+hBv+QuC26XVJ7/liiX0ILIOTuyL582FbPu8nlplnw4QQtK70SA3O47iC/1y5Dhu
V1c9OI3yMeoihrfOzz76aNH4l+kcMKEeOdfbFNRbZqMplg8bpS4uWuWgdP5KJY962xaxpI4NVeon
nlXKUynuNiSXg2FgeLyrjKXLEKP2qjc44K1MpL3b5DUSVFx/O5mG4gbJ+xoOAFh0eB2hLndoz57w
25toZObxzKv/QIyO+t9Rz0S0HBPI3b59Ivj3LkQmstPX3+wn1sYvLCrvDQarl4kRuVDXoEjqu44A
WG87jdCdXFvMlSfH2w9GLplgsmpxYogCPE02QZCCBzS7UL1oJxrPBl3Mx6y+Y2Z+3CC1fOPyYZTL
1K0o86IJtckf/lEa4TabbEGjMeZavpd5YklPYZFbslV9rh4QwNj+grD+q7VnTbHPafGrbM8kJIuG
hYfrFutyrYHO6MQU9BRA9gDWEj05grUGvtgxmbvKLIw7lOb9iKBsM2DfEP2DpIBHwOv+Ru5+FHic
7sSngiK3eYDfGtaMQUVwQsBlQnLdAeyCSAs9Md1Fm8DnvmvIwWvWjdhKdoO3WXO663mmY7SYszgM
Vii+dwBKE+Ey6QTU2XRlpl72i8C+VG2aO6TgPxKynjPlqoaTm90OvCzXyKwZeUS45W6vBUpn5ufj
2hlEE5xtxipAnTV+WFFrO8B38hbrRJ9S9caVqUSp33wqm2gM5lem3XLgI14XGSiKggPFOFNyLsIn
5MAVKeqiUjzqDNfrP3PGHujc7GP6Gorv0cv/0Vu8Dxivst80F2MWCcMOTS+zypqetPOFdWukflyD
l+OwUnihvijb3SDPnTlAZvCGFl1QlJZkq0tbV6fZznLWiiaEZZE/CdaWEafo7RmpU2ml3hfHkMks
f3j3jQsRu9FwPc2iHaKZrsKcwjB8spN3FTj841/unK+UOjxykeyXXoM70jdGb+TcUOkBJ4jE4A17
PFFzsRaHy+PMRtyUyIpOffvm86KuQvxZf8+ao8JZq9FZYTk/O5o1kSKGt6JSCmCGhUcE0S5v6T8z
ksc5QP3gPjlMEFqrzdBsklEBT7vb8jCz9fAz8xuMr/HI4E06bwuNViQVEC/7mJoNkIzeUkoYMZfK
+aCTlDvEjWRD9Iiq3Dbjt8cf1osRCdwgVT73VmE1XXpFl8tzBDJmYF6tLzQW4icsn6n9oxV8CQ2n
3ypx/I3dRuckj1ksk2KAABC+2WtTQpUEJCGT+Ryu4cLxt3lruGwEm9zcSgCDFFxCqX8XaIlSQGMh
26BRYbttL5tsus2ZAz/r68ygMr/dh3wILAlrqJMPycxGKvrvKeL3AiXwZLEp/9th2AeyoiDK8YJu
mgmqWyox7CZpakXOlpsNON8x7HA/nG51YRrbapXkbQJ4nIqKeeacEiDm0X/hEYKnhon/WmJiMBBD
PcrLQg93g0i+ff0rl/OoN77Y9gzc1l/zM6rNfyUagB7wMWNNXg3Tkx2agzz1EbLbIzfaFG98GUQq
nYf4S5gHqsZzNORiLqDaM2g8ElL+S9Gs8peuqtSQBlEXtKEAKlITjCo+7stpZzbri5HMIbGWvvFt
uaNLle+TylJUOAcWT64E6QIRGqXIYxvo6ol3dy4xgkh104z4EZ0mS9zkZRjKOPCPvkEEsw4xY0nN
bIT0PXT2gX1urQLDinRZwp7JRYQ6mA7iWnM+ywxUXEuDs/cw5c8GS7LoqcB/+GWmVmlDk3D/NDi1
W4imDAnhUmF6xPNujmZlI20jxJ6WuXLw1Y18uJm0SD/PS4fIJ7//LoLLC5znTOM3vpJYdmKv6/7s
/IhCZ0ncoJWCFHQTwym17NcP0OWgtYd1fp+StkGEnMO0gkkmmj9YVarvr9w4+V5FIopwRVt6pVfQ
P08lCPQJHkrzMLqcuob3QOU2X6fS/INmS0NbxXQRXyJzZlymNq0HOBIHowVH93TV5FPmfTpG1rdo
5cVUQMeOpMXxQ5a2tZYbJAsKguD5gQ8UMkg6an/HywuIhOpyBQoz4WlvCTTFgo0x+TxlV1VtuMXL
NgcXoj2reAVfOP1OLpUfmkB4xpT1z+GLIzNCC0IKWpe7XYqazyCNtBh6nxzgSy9lOEDyPKM8g9Lc
MjHCP2YIwZHMifJvfkvqdIiuXAdS0Mrbnjxjzj3u6sSz6Jkw8PB4cud4tdCjoZbToKMDxsSgbBaW
TxaIdrQXOYxlM0q1EM7FtKaL5VCdXXgNptK37DmaLWOwoC8GzX+B97H/G8vYvkDpcOj2E5806CS7
iC2tdwSDSZEeJRqByL18uOX6FuULlV1DDyf5IlKLy/T1vWz6+uv/2ZLu1JwFeH8DRIlyBQC1C0N5
Up0V3/b/nQasnzRyZV+SQ1fwnpZx2tBBr3F8KS3U8nDJO3VyxudYWuCjT+sJzUA50Z06DhDx14F/
vxHvFTnWlxpQC2idCFAS6tTzszM18cJZGuEsspXGOjZMjIudg6bbB4c7S9aocRFE7dhf1r6bH5De
ihj3XmJNudzMZuCSzattRaXFmOXX3r/25s4LfU6T3ZdyatnoLL5UiwpLbBz76b0Am4WjVzmoiVei
/SYGOqXKq/2Pk3pffLgc1Z8/jK5JJBgWkNDITGHB3ao83xqNx/xiENIM7I8Y3nLg96m+Q7LWLlcy
poAIK6l8hHXXQjbaC3odhcnHkQWvNq3+BVMkmEt/zaQTdNLlDx7zZtDH21rQi2vFXZ5LjZYtRJ8S
CsSxIgQ1tVGz6q2fIudznLbUUONklgrDTQlIxa+I0wdmB91iJhN64mzdZZcIcUrfdMMpMUA00bfp
LiKTIt5D3z005daUQPdndHlz4ewlue5KYANFTMtfGLrkPVNjjNJWB+q3RqgMa3gFjiGCC2JI23fB
uljNvFnQAbtV8gM2q7ACa/HGggzUswToJJYNXQfGyCbVl7mxnAy17OjBP3Eg6Hq/kuSrB5eXbR0z
P1JC5Vm90OJtAKz8Nz4/4kA5aC5d/3oEgtgAYemfJB+TLfAzeHGL+ODcBXQcw1KT9BmVJHZ7olT/
a+SpMb+NmG4SrlHJjRcXa0c/0G7kuGbxPWWfEG4Me4W7sGRD+NsGRFSgvO9CEVXs7wrAA6HBrOsP
7ZRWvpjZWdhp9SdguJQRKBlvfiT0F2GqwPhL+EX4CDtKBAGS03IVeSyQJpPpNm/dZWfAG3zsp4Jd
p9+4K7ixF52XPN/DfhzOzlwmNe/gEnkqYWKZrXixp6fg19PkdOo1Ky/qKyE4rueVSt1EmJ1k9plQ
UCq1ve2iaeDS70wFTKJ1VmXXrTCDwaZM7L+DQTeKWIX9aS5qzxeXG7KnYMYS7w2D23EQeHSKpJNG
x7mj7ZSrLST5GH3Rw2sg7hu/StHXK86u7J12QP+qpLSK0H1yXP2mtbJwVXVZhmEFhhTh7rpKPREM
wPE/oJ4DPkZS2WDoUoY+WIqriSh4ILIM8YwAoBckqRsUcKG4OD7z2sSztWvF3FA7UCLLVs8B+d8I
oG0San87sdsO9UDbxKv/6zCx3sYLXPUy2+TjZ52snEzDQZWRuxcHIoHRr16xLubmNCLL1W+IZN+U
sNbTkf08G7PxUAyLIveWbfSzZw09gdAY4SZSr4jfNNchbAJmf/kVYBhEkyZxEzjcfC3dlx/eZYiq
1qzjde3IUEHs2mZXDGdhhRV10s8c1vKZXebkbA/SzCJahgwsWHxQK0nhYUlH8PGo+5sOPCSWXusd
CQEGL4w2sRqyv/BntxO8Z9OfZMlEcjgWzS147r4neatoOdQGiLR7t42S4LnCbE7ZAT6HVZagBWqg
pPMrgTDPlf5U/D9Zm5ENHOkbunnOZQI1OcNTgrIbMCI8JLQXty1NHLhcQIZds8rViGilzPdP24mw
xzXiHPn40gOJkuofVA133XvW3mchoApEE8Sty55O9zjpDPzcVKhJu+lKfAH35kXrZ3tHYxz4Ibfg
7zdHiswNerlgo9vKtGsGCn548Fvo2wCluk8eaUZ/egJdP8dlPGwv9koRCzi8ql/WtGUcB1Pvv2jY
gLuxXUTlNKqmzH+9wm0M1HYpyUk09irCkfIIcUHMmYW/WkE+CV4BpQx7jVG2yLqedsKkmv0Hpifl
ANKURBJ5sLzddbCJKnRzhFzMpvfI35XU5ehiFz0m/z39jQrOgBLHQCbi+45ffTPe4BdEOqZQRVqU
ex7bkB7fXFcMrYI8DjSoEkQHCvUGyzdp9zl7MRXgV4DwWCX3LLrUq3UMnChdLT/kaPJkJGw0poX/
8dhpwYZrGpOVzwxcv93lPrxNhPnDmJ8rVWRaQERaz10x3nwc0USMCU53xl5gJLBFlXg2qGllKd9y
d2bBFW7TLdQBe2xealBMdbODHKJkvXCDBfF64V/vG669BtKnAX9dhRFepQPdkg3IWIS8RfIJMLIQ
d5dlsk2G9PulCO2hmiMsvG1i2NiQjNj+yfqpnqUW3NDUPFV8yqWzxhQWR3Ie5QEY/ANsXDR/DOHz
LkTKjpEwsOJ801jbKgNSwpXe3rWVBz3n6NwRdFwO6OG600WPfJ6L3kYAPywyVlt9emVJLkDRfJBV
vfhM+Lv3W0m7pD76sdnBfSpeRrrtwyuewPdj6Bt7wqDIWKf2jw89cDstap/H4uCoFr+FbOUVmVvO
7G8dUiRmgNFj0qyFMO4sxQgzT0LA9RuOOibUXct8tV6PQAzCn80SYVR69BzTiZpixT2aQaOsRjMj
1vjtNe/q3/kt3hN4Is36Iww2IH+BL0jgFoFDEGK7cZzJnviU8kB7XFIZObE8tvfRta+QnX+ofYfJ
H/ZQd1NNQnj5pTULLIeurbfocwwbWuGxDWiLdHLIfodDcUdXRnTZIEo4poLOA5gcmZ5NtPbXwR1R
3LdC7v9hxbm8asAeHym7bZV9wfoaLU75QltqscMq4Yu0QyHx7jVT5SXIyg4ZlQBN3585wdFF14NI
Rq+4E71D6i9gECsiizqQPf+CelbbTAeCHU79LP+yKnKwEZPwF9+glOatic0zeNOpMvxqezWuTMVz
7iD2KbEln6vOHtt7/G9PA8zk7vxYl7cvt5h2PW6Lyf3tYOcW36Klz8yDNujmu+tlbtFednJZL9ff
L6Co8r3ZCkSiKs2cDuqDey//fepZ2iboEGXFvbxNQWuyFSqVZxqSG3x24qoBRZ1ly8K9z9JcOL6f
bGn+KdExMtSRzUJzCCW6/LYrjkRLQ69lOJyPyQQr2gdatRiVS3ClvaQWkAhKnYxVFCQyOv2doId8
UI6PXpe2sjCPcJBbBFoScsWZn/n1EeTseErSGxmyLMvgtIHdIhkom6q6wb+K3sUTP5KGCFhUcrdk
DKAWQvOa8DDdISrQyogBgIx//rdNqT5W5b2JvBSRVolX+b+rfcqHXC3ov+lWAEpFLLHdB4KvWERX
/ialQTtn/04GZeRJYIJngBujuuREJd+BwVLmOTjjOeVNy3jKU4ON3BNld376VFGJKkF+W0lrJMrI
14MU94Ar8KCc5nBqPb6SB/gqVmDq5Ye+71ZA9nmD8Uucy/EJdaPMMu4Q42OJMCYUlGmRRrunBZST
/hpzWqtxEmjDIRGbfQ5YWQOnbdkh7PIf6q5p3SPZpV00MWhgcSYiW56NmIAiLR5E4Xflrew9D9Ld
DlRXWo7izMLYWWi7kH0/TJScWIvE3wM595hjKwb+d785B3kMiqYBWq+A2FJ0aT78cjSxzKAtUePe
lU+auqZo9qFhXMNp/v9s296h/svKBCD8YF98aZWP4hRzdhIRbfBn9vbAIpAHCkCuCIViQZ6mXQ1x
mGvyHnpz/nrk+l5J5YXo88xEM//sGQU/Q2Q2wRmq1lgI6Tk6Yth1hTQCXSI0lK43OABYK2z/mp3w
CZExYWdfBDcZXFhsxOhEMYHA+3yekBrb7I1wGoiEF4yCAld/BDo6XVa6PSwK71RdSVRZtj23a0mN
XiD8N55LIpIUNk8THzkIJWopzQhlG1zS3M0QHYpreE3VqO2rblKon9kriBgf/TfsA4yy6KuJiUGa
VQpZrVvFccPf/pjAjIWQTjaHim8fryrSmFtB5uS1B9bbUlrANmd13OevOizdHIiUJUv7HklGuP+k
L+L+Iu5I8D/4LyDx218s99HDKAO9Tq+sNxgYuyPM2/M0HiGin+UM5hPRNtYf1s+DqvYTB64QtplJ
C+ZCy3EU9CddbS6BBaLBsyvSdj1opt198jAF/NJ97G5Xq+CFUzbobtK8PGsJqu5ZBwBpnNF4fRUH
46QHuaYW9QMvcl+B1SupvfFsnl0m/vqW/H/SlDRN8iDeT6P6DooPymKHorRmlmzj0+jkCI0FLN7E
qX88xuYufeB19Go1REEE/JOS67oZsyxid9PXhtAgRZPI9unfiCSIG2MCFqipVajlAGiyLREnFQE5
Prpq6VHRQONvi2RM9zcaeLjyfFOeTlGdBSv1ihP9V1NVSp9vBDzZ1/0Ds0LEZ1kEl5cqPxKeJnE9
WRtzXO1YAU0yfp8F7uOX5ArarPntr03E/RTP7AStG1WuWlaySR1brDbEoCtmFKgObFo8IaQ1Sp6g
TIKzzqXKmWYT4zlGarxk0ctbf+9rt7QMpsQOpFplczNVCzTU+0AO0oBrAVRbzvFQN0OF2fKh3rO7
WIzo3VwhABcm3kCS5gm/YclpKNhleQuh3XhQISbNZ8CLL3pH266aNExjyCOwKI6cokBkjzsoBo2w
Mgpv19+Aaa1Yl+o0teO1DFsNOPoD1KlyXYXXyFtQtYKgOjxc18t3WwaMQHuVSl4ESZsKfTJ3OdSC
cS4wNQyi1juY6BCoMer3j4TdgvkSWCMnDU+ARGBfLfSrX1gVp7+C/OXJgti4Sbs0h04jw84FC+xe
6bSKKg0zh2e6OZIQ+LWRzyRFdeSbso0MWWSqoNx0nPAleGlkbNrbuYaSHVInqrkk0QXSkOTaniB1
NwIzVW9jFwgPZgSIt5pSyolsEGV3fCMelv9ZNwLVcOmH9ehCGshIyonmlQPnSHJeT19sZotiHf1H
o6Ni1Sjcs2V/X8ffrZyi9mbrWSzXc5ldsUSzvuUL7YQvI1KJD3uYwHN0Jimlcb3Dt5vV2Vpn+IeJ
vuN5VaniZoLJn4ohyFovitRs7ER05/dvQXUeK1ISOUJOnRlGnyOdRXBTb7MlhXEF13ZqFURZCTjQ
pcLbeIPB5anf0q0bjjlUzoq01Dl38mIbWKkCykquFU9hjEt/kugqBfHUxa/naY+CSTezTzTZU4hs
SCy3TIETqtFPVtBYR/04VrUBAczzKrscwn9WzDNUnJv+XdbWxLtNxxu5fpKv9MxyBBA6sOeLqk6J
40xbahvYK3ipDY3/6RqfGyM0gVv5stvGWpt8bKf3k0sa68YL2Fz/aHVoL7qZaeYZuv7YV2hKZ4FM
F84wjOSMkNB2A+nSnTTRX51qKwJpYN7vf9XRvQpRIhw7q7/koqd3CLZD+X6lOT+KvnVO+qso0rOO
6IuRYLDKkCGkq9MVJ4oN3Uv6q2afrdLySD6f2InHpnZdKxVyJ9SGaKrd09nVCy1K3ghvWGmHdxtm
JprWFyFcQtAoP0Is52RS4KOQ0nUnBV8wCtGYC71F6BHTjFBs1n0wyAPQHvmXn1xzi3J1/D069as4
ZYvXIjHLMRIlx7TFkBJ94TehPgEWEnhCct5aQDYxhIegCa2KXS67/vZ5r44ARi0hyhqu6NeSWzwZ
FcPQV7v60EbimzSp2ttKftqx9wVZGipvyo5QOe/05Wn+NNueG/pp3Ri+cBp9ZXTRP+DrcRhYCcNq
duWyGqn1oRaL8XqIRKeg87mOZZSpDEsAjEZpo/MKRZH9koAssYoFmeY0hF5ahPE7iVpVbAc1yQ4S
/9H6d1FN3UB1Lt32Cw3wD9Jgg/T//GYW+Iw7v1FFzsbjrgf8gw50KRRAYktJQv8z5IUI+7fYUzNY
nSctVEqD12x42zAARBtmWbEe6JS6znEV5YUXSBMcxXeZkP9eBCs7UOp7FKBvh8mCmXXH1VKBuddt
LMOSsfLltKtIf2VDK1zw6I5PerxonQzLPcCGPygO/B8DIga6IsfINK1e07wuQXWbaeeyWULOzJde
1t3fP8FfVXANW904+Cf7/Jg/ezSOk9/O0gwFxXfpQm/0U0gUVTGPbREjz1aWlZNBPYj8N6hWOmYl
7Nx6r2kj7g4AnhW2O8WArFW4uGGFDtdeSIRFqL4f/yTDQNt7fUFp5i/ZBBUfEbq2YKZllLL3NkWi
HPeWfvLEYlLylP8q4j2uvNpNAIz1bzCioeJECiNgP190dQvujedr3UKcSYWLgQy9YgYZlr9VA/ui
MWwHsb6RWln/jGQrJh479fndz/Op2hSrg1w6H/hDRBzpn27MsKWwvmgxleSw3e2rSO9CTbW/ZxRH
u+VsP6Aj/yo5+9dwSF9y3xlumk4FDozO8Y0ON5gtMqeTkTbtUYUg9DpV+t6vVVrUhX9i5Yl288jc
JumBZQ8JNfY5NB1lGo/yX9W8PuJqDoFduh4y8dAh1c8kweCKX6yfz4nSQsZAlFtyS0K6ZBGYZ98l
0Wec+UbihlzM3qliM1yX1ldwoRCPfwrtrBS8unzBT0Du5Po6+/kyPBxffj8cKIXELFnRm3F4gArU
RWefE4iOjGCZp8BZIa2YUTI+f9txQO5yI9kxPnxRR8Qt0bFrxBoZjhthJ8scK2NQWcICwaT7LXz7
Sa+cJLUg2QM6JPUPQsAqA+hNWKGGEW7X8DBtLM1g9I39o7/lhhXADZ6W8WbWfnys9w8SB2y9sM9b
aqQy75LNObHxATZyX8mID4mBD/Kk8K/joczqOqkErAR0QYyHLO0SX75Klh2b5P81NQJb8AO0ocki
5Y1pfjoxQmDfa4LVeukLtfU6ljh4BQb5V2911R8Fo4ymD5qKn3Yso9AXXJ3jdi5XgZ8sFsxNOhmS
1mSTRXFdtY4qFSmaUXBQ1gIOg4s5RXlWl7s4uDYwUuQ2YK5e9oCg3ngGDBjXApvJBYUL3xvRqxLo
giRjU7uefdWAAW7RgpAt3B58y+Gl842sNDapUFts1u/xFehwiZtT6yCjmk5cHBRkO2eYZJ/yDJiQ
YnYFaBICQQ2B9/PJpRALcB94+iI1uKVT2rEk1rX6dUqcQvPdRAJo0qFUXkmW6ZBfzYQcRchaLZYb
5AoMVlJXEFzNPJXG27WZp+NAAGwTIvy3XVN4w6MmeDJQclfBOD3+XxnboBm1+ZgZ5t+cH3WFC94C
76XIol1ApEm3cEr9FGLJdmDFqHazN7iPi654ql8/dQtlNipYfmRU2uzv7hA+3wNSxLxycqpwOXwC
W7Q1JfklIIAg+yx6hjj/RfOblGQBhyrE8qxos+GWv/5aiajhGdumP0oahpJHrAiFnrZO8Zg8sSzR
k2KfZ2H1Gpyhzif667XQRyftEXJVujIMCo90hJP+PIDoQ9QacVcOQRs53NhotNoa1SCgrYmNd6VJ
pR8Cafw9VkndXcJkNk1V4nZoA9mGxk8ZsPyoo8HfmGT66dquW3YApxppIYqiU9KDDYAxf4p+SenN
g7orA/TfCP31JTiZJhHUFWSBZc6niRFD0iujQ8ou2V6sgODZXC9EHaJB64aNoYZfUTnYLfvC9cTw
BOJeJA7ERaOJQI5Nl9BlaK32DYy7szJDaKwVh2oALiNUga/JAhG9XOCeY//v+mM7IZzUGOzC/j9e
aSiUWsEzX9nDmXWJH6SMg4yC3CSYUjq6lTYJfsfkEI8ibV5mbAkJlW8Qjm3CjTbZjPwecNNo+/WX
lWwVpfKwNfmEJRalTavTQ9Rt9wt7NUFPWplVhKh3Yc6f25ghpwYRraotv7kfPrAHuZriR7qGPnKt
1BY5xEFas2AuOm6OwpUuqEd7IkF7F2b594YguqhoGPxA6eyf6tB/nG0Ypf7lMjEXZ8e7Pl/EWbT0
8g7mjpe5sbmsBuPPo53TFWE12XbPpQhpISzsyC9am5ky0c0sv7T/zjzu/fPLOal9185MKjGZqhkK
Zy8O58MxIroK3nT+DmwrUzKXSuA9Afn7IYWZxSxO52nY67i5eVVQRhOLy5iX4w5DuGqbMQCW5EZP
Mgk1sMpme1bVxZaQ/ym8dtcnr3ruYk2Kgjqo/y8ahvQgih8B3kkCVsuhCLCEVu8bolVBdfbJg4Zx
gxed5MRtVzvnW/zEE/i63Bwj4EzqOu0fqxOW16ozZ5ByjssaBdrlKZjRhOxjpWsIc86razip2f1t
1aqvAFAQ5r7MI5oYBuc+73CrNKuAhu6qS0luX2hZdPhorDpUixj5NQ2zqA7Uj+hckXxSkkIkKvYd
jfnDSDr2L5wZhTxXtNH+S9LZysgOSMqm+12qq0ESFw7vHA9aNMZf4KS8mMX3N5VlnW4AsGGDs8+6
42/iceGbhg0tHZ8bUWaKj9Bvs8+QVh36UYPDUDPa7ouvGsWdSOd6dbCoTI8RnhZTVK4bxCcRUesM
6C00jt6y4T0XHr5upqdUEX7JUPbNhLkBQEFR+OZkGLol/M/lgYsaCYq3E9L19+4II6M5T7Q2gRuU
wQJSvaU7sqhq/EAz+G6jVn0XG4YSNM+avzkL4nrchhLuoTLB4tYs0ZxhkmjHQHr+JmED0NJhBrD0
xiVSWvUJT5igjAuLzyzO//IXxRk2E5D/KXkuDzZ2cdg2t16ItbboCpiRVKay1W0bbMfSV151kSk5
VqVMhxqbQ+K2etTRaIbRotYMV9S92B+IiNECOy70yqzszKnoc2zYy1dvTpJQCdHUYNlZm6JJBfPd
sLYIxrNyk2/M1Uu6fkynkRmxGrd2FIrgIxIzM5fJoifkmOWMUGkHvQmFN4yhZM2RdYfSbsj0Ewe/
Nd+Rnag7K4tmdZ4XboHV4yMmGZFgF6Fof6k+zOCqyFOnJyTCexxO798/9yimenPmQuSGYFV+m0mO
T9xQDlWBE/hCdLZv6lkxU/jo90VhN8j9PIp3uy1SyIhPhFdzw92jeN46b1vYu9x5gQJWL1aJCiQ4
kQUeDzHtx8IFXCMZtAzg2DaaeEkoCxnIRAxPRIt6wm8oEwVJon/0DERCDfdN+lR306ntpdx3Ad55
bdLAZgmvOvPyjAxZnLISp9u6QhEplVtLAjMBGCg/edQptLuI52CZ54DsVmx19GL4/aTt9VPZ7iBv
AV7QuCz7QXcUKPxwswYaCsQVvOgpvJl+Hq5AviE5X+BW7um6epyZB6otJ90edKVdr38DkywyHVBT
NOn5ch39qVn+4+/nssGj6zNxmf/D9jiYsEKj1yQC7JEb19G15UDYZ4FTm6mRAR+5U9G8mWOg2o97
9M+A2C2x2Z4Ol9kzzr2ShhYE7T/BDOf0D8ifTVDfdiltgRmDkZ3jGY3c9phwVPufTC19eTcPbHii
Xz7wwB45adivahTQOW/Bfa7Skm20Zl+rjbf334X8PxoKeQF12LMeYWLRXTMGCkZcRwWB3nfHhfN7
v3WqQKyQm28MxI/iUR+u9eYUxf6DeBpHnWnt1jIeuVyG9ppA6bL7CBaApf2Sr9b29uq5z48TE5OM
W2rV3CmAGkPAY9es+BxCweBIJ1QDqWcxmB5HJWsSIMjaQxGLqIKUyOdi85sHDI3zPVMdw6ahViyF
+nTPCEKiB5CpziXJXdVTQDQaN3P3XJK0ydpC8Pge+ln1IuO1A0kSO7kiGD7ZzmGb0B6GzyqW6pZi
dFbCpDAs+By3xRxgHdt4vZQVoNE5G716Q+lvq7Xz9MuFZQMTfW69r9OMcf+YHTxAhKCCD8z52NRI
IrqHGI3is+UIJqfHsEuM1hLsZg9HZxHwQvDgjVwgcf+gRHo1/+80t+cIZr++gGcsUvD94omEXQVH
t0qSjwhBBa8/36FkGO7PWsZ5ylAanzPTyKuKCEjGCpOyD4aoI5EuklXuhrJbIdcYFl1tKnRsJtKu
MXk/SJ7lPUSM3UtPW7l+SH7/8muITlgYSVGp1VyF/2AzNz59hrwMddmai431xQLkaFr0VniBYcTp
hveTBxc8YQ2/O/7P+Pq/xLRuC4y8IePPr8aUs1+FTf6s4xpOk4g0tMT519CZZqg53aygT1s2ux34
gRWVO7h3MwV3sT3pbqcVir+kOMh0oADawCvAmE2DWl1AURflPaowtW0xvOqfnyE0VtPuyo6JkfyO
vsaYUlwR/VAtW/jhtM17rNkgTuECTFCUiZcuR6MdfjUYXpYsUp8SCYgLnrqOREfjqQYCmZoU9U07
BFSt4ZRYgf403spYvm91Vv+4UwqKA3UMSb6Pd+6k8MykCEKNCwoV6npCT4M4MBdA6fxXIuNBpY5l
SH1APeSYm7fBXWLPzFhi9jCVLFP1SZNaaboVUp6hmVIIfx9K+mse3HH5M3ieWAlIxO8RulI8sivt
N1q3Z0T73tcO+UJlBIl6zFqC09OXRILhucHf7dRjy4S6n1TVFijWfwo8mousJt7rbJF309pUQp9H
rsaoICu9ExIvErEfuUAHuQ4kBWnWfKH2S/j2z6GQxVd7aCeQRyZMv8qOPodOjycZNqYmYL8ahtSb
JdwzR80ejldR07H1ZHsHLt/fNurLLtzeAmAVWjU6VUeJnieT8kvCwkXgLeBwDzGYwnvpakLevYEh
a6E2g3dpWSK3S44nO9sBMVInmDvUlVNusBNuBR2tKiSKWrcIrqCg1yXCQb/qbWJsPF06DhwP6ZwM
gUJJz+DOGObrLIcmnVYCvw+tW9ZO71qOo+UiUCmpCYai58B4C4Z65ccfYfaULmKbQ4Ch+qjLIHaC
FDVg7m/5ehPfkGEZznCZwhORMM8tXB6W6TQwVLC3od9G/s8Sk9h15AerJ6w2tPWEWMuTyrsxNLbF
h3IFlctoQBs/7DEMDt89ZDfqUHan35MNssgUQvWYArF7wlKN3VM7ZsDnvmQpOavb7P8npvwBvdWy
lGv0EFcWbHk14XyBj9RRgwjcwC9EOGiO+4vTKVP2F6Yekjrbb0Qp75wK5l2MBWtJQQxJehWPPgMx
+kixgGmppQVvUzzx+9zfL3vIjF6+DlJKBdTyBgBUawQf4KHXxLufiu5t4DoVz3wp0EnBiR9olqLL
9Bp/47HJBL91Jcv3JZWp4IF2LDK8L4uYxyW/WJDymLMdyWPJnzilBFRdEj39RRVKgjSl0Nf8Rh0K
FTu2+N2TA0MqQ7UcHOh+zyUnRMh3nW82yL7cdKt1r6b04Qn2npAk0v9lT5DDGu4rllvB3sNep7J+
8ZpRr0ZAAIY1ypPBa8qcWfqrQbYYuO3AZa/pfVLL8kUKlU68ER2AP9WbLI+jkcG0vBtYN8UGbAMa
zFtRF0C2ZAZMnqZ6oy+WRevZ3zFJTZouWOw248hiB/CLCH8Ml3/9i8BBkNZOv1Yqx1N/1IjnZ8B2
xbntl1qeIWN0kHXYZbuc7/HsHY/VXpSrogTslNyrdq/gSnCRthbuayUkxhthM0Hb081TWL5YT3gf
Deju6cq6MNCdNkBKhWbkVM28tITvVBpLsEQIHzgrqwwISCnbh6RgH+CQxmnxE10roVw93v9bFpyG
nX0wikuhITo8BhAPk2F/yUgOLKhKex7Jnlv12iDAjnTslneyn0rxX+V7uyHHN7x3Hd7qSw9QCrfA
zWfIVO9le+kCpJhnbiAseTNT0fNAEyPOnmOW+x0AQtCvkvY0E7nswNqdWQDcyqu6DFUFmntgWh5X
qnyA8JjPq+K3rD5ZnCDR/RaRnv2mm99O3O3PRA6vk7CQcigAMMAycS3h98UDWjGPbxX4gmNiEblO
QHJhr88vjHxI1/WAkwxc2nCew7JaBWz0E60QyxSZf5jEbATMS94DlFKBwk0ogaMGJtmzFy9Onnsm
qZyuT1ikApeb3XMZtx8dOOUXvKAT6JpLl+jg26ZDB/FGTTnI+blekxUtwk68ChOxp+6n1PJAoqpc
fNLiBkId3/3bhyAogFTrCTQAfV3g7EmsL4ewSNIZlHPG6saVZydBOHp3nBKee5W2wPkR1iQpQdft
O6kkafEmGTUXQLrzLqpP6ODHB5yk7LkEVf3Q5Uxj4qjOhkqtlQTCSf+s0p5tNaeKFkIXWzJxqwme
zbIaGP44CwBbMzk6jBYCYCznsffME8KT8P/JpWvEgiyBq3K42HSdwQ/mAs2qorUfw0D25dFbwwpP
RtjcpCWyp+rdN5ykpdElHNIOy2BVvnUgEeWjTV+8mR9qgCsKGZStaLGWV0VWpQal6lDd7egca6Fx
O7YITqctKD2eD00P8Ufp8XL+NxKhCqxbwjmEutnKIApIUtBhTvs0mjGj+3OtVLWzBflSP3JIVZpL
naiBaatv5vIRsFGEyhqnYqQmsNqLaWgv4/7kbTrjOxesTz20x9Ohu+Som0rdEkk2A0kI0Us4JXS4
E07G8ZZqOZsLNZDcFTVkC/YkqyqlJ+V3AzhWLtA6tGHwdfSKuWvR5Fopaoe9X315hQfXaDbMPxzX
QnbWHiAJ+qHer4+k/XowD0WsFqTIgoGAKNi9Vvco6MftsX6tnujfG1EarynQZ43iW+SxjNJrbSea
2Ffgz11kwuWrUGsRFHKQzGztFDz/fdWWiHqgSHsv92GTsEFcOqCYLtVouQPDVjVI5gGnP+A3btU9
XPzMKSM6E4UeYNCVwJ8ku4EaYxRILg+ZDiSGxVCYipgWgqbuRC6JKIEots5vGBHCSXJ1iCO8gggC
NsmwL6MFwt0QBYA2Yzcx9uJwjnlsTxrzy7re5+gcohh/djsl5kx07uwKw7ioO/IuyAFskWzK/2qs
YVuWs5qu/VRhjtx1HWjHXL1jyLj1d7nU3lOU+8r4yBrA5KLCNKCQOfYgOWl5NfyhPKGVIWB5qzFu
WNg/HgjUUHvAasEHbJ2Ru6L/tBlEbSGM0DMn4OkClV1Q9fLyPbK4qHXsjEa3jMR78fuSYbm4N5Ed
u4cZIZt4pTaqfHYiqMZl9jI0phDHFPomxgY1P62zVU3sIibErBQCoIpUoSQ8uBM7cas/aqRthiPx
B1sT9AHZ3CpZ/NxGiKf0aAhkJztReFb5O0sDq01IbxAcQr0pf2wmF0YFafcFuU8GXS1N46g3ebbX
NJaMcLFd5xt+rrKhrBmmPTdWqOC6nmwIhGxrqcTPHr5SUxQw9qEZWGerfqjFKy3YGz0JVMo90A9P
8dmYqlXl84W4PiEtwwHF7t/2/QCMcgAo8aHJqcRXWRTZbaplHcbJSZYa3z2I5/L2wDCV8UdAHf6e
EzN9an0u1w6DN8eqS6yS2/QbGBluMPZDWxAK4mwt722DaT2pdx9E+v39usqIVC3Ket8G0xDfTc1C
fsfLpvcwECqSZ+MDi50+pkPeHUvIArrnFfIfFykDh/jLLtUu71y4zSpy6wO32wIzSNje1Zhqt37M
91bkaODSEg0OKjkWetgTSjKIi/PVu/WyuNnja0dA8jchJZDVdYXZph58GOear9zRLtaN0OkE+FUd
XK95iHYQgJPUGVOIrNm9o25znIuOF7TafkEiUo9k6etSCCnaVAUJ2Qrnsbc1uIikCGAZ7autKzKj
aZvuKoSavIAkHgsnjwdnKbB1B59/0yKeJInijHBodxoF2kI8JLljMKRySF0rvqnoyd149H8vq15A
DhCuPvEujcwEG1YE1Tho9v1NzogYMhu8o2zu6+WIiBh+Q1zGOUBhk993snFWPSw6qajnDPEZ8igX
FQQkbloJfWr5Jvn17F+YlptITx+aUiO6RxwMwecaPu2l4mi5tR4pXXnmft4iAtiWFxdQBqZjS7Kh
DwbZfUwWg/BhlQWJPsQFtYKzPXqgWh+Pfoxmw6J8jfZiFVbiQpQGb6d1ZwQTUWJr/+2PBbgTUYde
VoLE8rovc2RbXG0+8uCxA8w2HbFKMWKA+OJsiaJzsgGX7D9Bi2zZpF/spschvPpz4/9tSyFh/MTr
D7rAzXvnYRn9qz8XDzaW/pYXvcjctJueIWm7bL+nD58J6V3xAWRSH7QD2GaKGqNWF3ZRgtauLnMZ
UWNYvnEyDudc7KEfhjJqDYo8iQ8YeP7FAReCgTmtN07n2MkJ6QSgAgCqHZ1SOKVfBYSjEbNyl4xz
dpwso0vGLbz7YEv5dYRJ0ncR3WpYVTbqIxBepj0YehRB9LY+vqyxhCOMsJILAmqwwMwXYxNmq+dy
tRV8oJrZDcGdxq3J8IXdhIjjx9Nla72nmMJwePdF5iv5gV4kN2XMVrVgCx8YWnusdCbOZijoW/JU
VLz78Z9ThJ1BLsIxalpmo8/hCaGCH9hmWGmhMZPwKk4M0zaUuCpb0521nWIMcKfRlM6NAIBd1m5T
Mtd/Vpx4BS8I4KhoMdmtwEVbBoJMnUBxjRp5abwi7y6MPqiCZcsjyuuTOGCa0luOuMFkQ8aB82q4
NfaTHrbMFSkx1AdNvsdeYDbZDbSHA5ccYHyo5ZILd8QBDTVohUL2oe/qqpedfRfTC/azQaKi7SUW
OAPFfyzs0TPfG68SzBEc9cW2PgJT9IyOClalz0FnGrpWSgu6OlieVDhjhBDJgSn9ShxWIIDiDN58
VbFax+6DG86Z3VYd4EFZSYFKOC8pe8GWFRhrmnjrjkU5WvRX8Wom4NOfwTGLtCb8IEbcxNY8EHQH
X9Pg40L3mdMb/6buzWaX/Gt7yZoR/AYGbhgmEVmYq83velZHI9iV69yQh/mfOO/zqSJ4sz574I+I
9DGg6dZi8XuZio8U+0xh8jQh0QnQNUrwkBB/tpknPNz42DPbWrX+WtaTqtprY/SQpvumY2i9hbsl
jzVbDKMCHscSEJguhnYTDgqHomOKwQoKmB0lHfvCj7YamAmS8ANWnjonDuEMkep96cayestuJCAD
9dQDz31mlhICOmBzyv7OvXYuqE2rKUzi6+qQAeJqE9uQ3dpf9fP22HoQuK6tI5jHqLrjGQfgtnM+
+iEzOdcQ4vxlp8/6Zx0Be/a/CYsikjT/56c/cRSpIlmh2cHmW4ppnZyKfxGP9ynHz0Pzh4gbK01r
6JhiU+SSMDfhK7zn4l7CwFfyFFL/qBBU+pzib+QbiUFrj2oLly1A5sfy+ne2quibnZ+Q4v5ikkUY
cJQvVuZ/4m0BiC3AVAcbkvhkrq9E3V+MN3KctZ4NFKEdoRn3IfXN/6eB7LtR1Hae01kxQN+/PDQ+
q5part97fKdBtVacfzBtkWu4RtipDwj8PmUyKfmrXEtq8CjTO6h+MoY/g2FMv+XF6jvwV2mcqFjS
uBjRPSKiZq3D6gHWq8ytT1KBYtIJCl9LgkCX4AjvjzaPnYtGodcnDrUBmNAuj69+24ahvmosK8JT
mkjLlpTliDI9Hg8ZpaOmhbtLcYvIA0b+w3BOUH6uszZrx7/bnHAdS5cRWaZZS0gC+UaSZhDc3B8s
zIc7T6SLjCLKGGJrHrjNx6MUbvSMARPtet40j3tKdWeDQ1OYMcfCv/Jx5jdxF/pxFK/77LWB/6Pg
T8ZjQN5iAr3X9iuNiQQyA588rAfloKixnHXoU+zQ9Jj3tlo5UwPVb0/EEDY/3+Dt96BN9CJrd2Od
jbq3LSJ6ZSR/uKr08NSNfBHu2jB/QNzuIztH3WFAFdtB0fv7BgOtlDrCnRZqb9ojvvTZS+VCcteB
6IJfsGFciOR3aW5MVhygKIGrpRc1vTev83j4ccjr3YJJvbnz8g6qKvLApNTFSyTyh+mhxJpalmpb
6Y93Wr1aZM9j8a/AnWYSMYxAh8cgt40r4pFtTR6gVwiHkqn0yG/A5Z+KFIAoB+Bcq8TiK8EoxT3j
4OJQUItY+qXv4nRMeAoFIOUhgv+IF9aGLG32s6frB5ukUbhDZpD/9iW58xvI/RfBWYW0zQcswMCR
mhGT3B8c/E1DlI4/pRbBfQb/R/nHH/N0ZSzbkuqxvuGGqYF+4ijwzjFgypyLUQrtM6jbIuLJ6eQT
lKvorBDuFRQC8Ts8QbLe4aSseyuwR1/XEXOIE0Fe5Dx8zIOLsmzFWPOvLwWxqHAFC2lMrQ7U5QXV
h1mkAlI1ai8MJVorwOQYjialF9CgJACDDyLFU6LNxERtAY+knxoLSkJo6SptpMGuylxVAUjb4wSt
9OV6m99kyZNHoQR7rKih2nPGAL+tqWntfuDdUWwX707a+EQlZSUHxhkPz4V9Neu6+mzblffKK7B9
L5QPjq89g28aiF+5V04uW8DtKV4IaXyYa8bQLiF3Jvazu/Rc7M4jyH2KE32Kc67UbWFU7AWAdV7p
i7SabvMoGzBmg/fNk3r9E0cYxGDFHDU1GEvh3A+ZZhi6Z7nLTke8nvhgXlhb47lWgmk4IMQFrCP4
Xlrf+k5tp1mRaIkx7Jqq0zBDA3q5RDWrQHox4dZyzJvmGxJhOxz/BTfZvPwW47hdfuNoxWM1hG4D
5NJeOnu9nWZUO76PZNTVFGnT4zRzV1Da1D/qT+C9YVI2VD86H98oVjo9SgKdNWMRHx7j/ObAh+8c
Bcq52nmnypT41qkVxidMIAbizlUuo6bw2UtgqqOPvwcMyDXGKuY5IxyzX1j07vpdZ/nLr8WjDhVX
1u5zxouCuKaqeWj/rDd9hiM00wiEgyWX1UO/PcljxOB0JBOK6Jel5lx2esMZxA1RBP9X5ge9NwCJ
nIu0yLq55h3uKn6tvsE/hs5gZ3BunbsHm+iEf52WME8TsfrGR6SAM7R7vIczOUADQgzRf1E8eQcA
MELD5dtMeEREi8rbNTcP2U+elM9aVcx1M5z8mTzd8yCfhg0NzwdognctExU6ao6RtvNSKlG9WzEf
QFtjnpCw8Kcta+IT4xOpZgKP5JV/j7sW536tPh9RaJzZbz+CwwX54KoK0iu6f8nQ60zsvQrJchKm
tTGqjQ/tB60C1LbFCUhN4xe+OSpK45M8HKHRsYRBfD7Kc8f7dTbKtiPozQXILarU2yFeVr7rTKoR
jq/OG3vSgJ6O4VVCDKkuAwR5dYnbs2oE/X9UAY+QVFukVfmoSnyS9v3+RCzlLDz96eV1aWkWOZP3
yy52UkD5PlTnonfOhXirKJmuOtYNoNdfJz2cKReQ3I51EYEiOG/IjcbaTi+svgttlskl/pxv1zvf
R5BPOneZi4Bou0jflFNZJtLYTL0BTpPBY3IRv/xi+vREiW7GQAi3v/VzwVAg9wyVVcSrPsuNIR0w
tDAKK4ue572sqIiaLEEqvnHKGeDBdpOIkE+OCs3NGsoW9/64lo0X/x1CR4toPN+NzwUIAo8LcNv5
lcDUgyhqx0xNWbix6rNAZyVTgLGYBD63we/Ng61nRGy228xt0aTjPl4uXKRFxkT2izzBjWERpvWK
P+2iIl7pxCQ4LxT60z476wbMPnfGxTSsqk1v6GIH/WBm6tFXT/nqQqekfPJmlbe+HvZdbvrWhPRs
RjWkNuW0GjOzBDc+DAum/oL98z/fkHzmbzXi1j8S09fPz7qaYYFhVBI5uHh1eLTZm4vX/xSKbVQt
Jpkl78npnQuFJ2lbeFCmelIhFrFhv1gV+GrQxzNeV7C+cHiPOMTY3nbLFxpUME+bnpzngv9ssa9k
glj2uqKs2Rvuh8X1ZJ4znJGX9x/ZTsMoI5YaKIdF2IpUHqDesXmS9TbRJRDbLWtH89P2rx/jifVc
vTmxuWk9+WJBYLnmY3BJYZ8CEGQuTfoe5hXwHrUbRUNCwOUg8R+ROPvPlO92HM2LcPKCkrBn5spi
SOpwaJ/XKNFgtMOK9bf0+A0q+msswi8hPSTks3IlwmdZH05u1GGr+l9C9LtKtVHYxiq1AbGxsS2a
sB2UQlS60wZ7cZgu0BTSNV0SGikUGiiWj3zzbu4JdIdRx4/5JB+4+SVcxpPhmXKBjDukXXu+KkGM
hpiuplhWI9vI78e4NSDchm3FVb+/Rce1vTGyYp2nRR0pCJdPUux4DkXBjVg1+NtUaG5w8HGpOMpJ
dO/cyIjYkDQHzLjCD+ouU/4e0vkfHnJOtZylbvAZGdcUnFoRA09tgI18TrQq4WW5nCP9Wov0azz3
eBXkb8xE/6WYj8la9UISzEN2Al+lw9EzuqXWRxNNHC8Q2yD2CA1FNT78AUJtpDLDjYDsc4GRmGiR
Atm2HeEcIV4W5EDPJiqkQ5Zh8yEbnhOC/Xg+VAmu2tRhooRjVjv+wY1Eag8CT8G9ouGq3tQSzXNq
G6AavVCbfj2p8dxuAlPUGYiktNnUvJ2y/Ii8Yh4KDnQsLXxcqZr35f/XkStc8zkkSszWHLJAczRV
Dsi/p4CxkANWAqVlyz8WkWMzpLNgf2BVQpIAsbZlhF0Umhfbah9gmvCEwypcnymcdTc0eoxbLKsh
0oxXN5Jm2DE2YDJFawMmL2JNvpuMXgsUTY9fbErsF9wKNCh+GHC/24y8Gfu2blBDm/bMkX3ix8K9
OJXSO/QfSPQW39I/DHH4WEA25OEt0zw1fIkoJzrqM10ZItnRiU8OOFSl0tH7NHhzj6iTQqCosbAm
p+zrfmhvoltQycgdVRUmcOQ42HAc8PD5HWO6KOy6d5saSNCz82z4HmF2EtR3LTdqC0e4q88mEtkd
E/QG4yVaKhsfm5BVht89VqTzne8DLZTj4UqW2qyxuenchXvRFbUkg8BISAl3MqGXUZksdv2GZTkU
yUtbQs65+v0WjB0fq9rLoV1eSbHz1zafE6HOV3cUMdi8B3DvEKCNNQNcuz8vY/HPPPrwf7AH9E2h
TEAMfB+xxO6Yvtsbidd9CHCAIDeqA7pXPmBh0MXPiBu/0y1XFi79zIZd4jGv+ezaGTzE99VCGTsA
d+VNEE+JOIfQBaeoAQr+Z3mErgm5ul8ygMPgVman8b9HVNtHLIUO6O63T2XEEx5BUdwQ1WMbMqCa
GsbVsLW17/DuVlyAHnRs5I7/m/f5WH6sXan4H6lCwFD0Wx5hxSFMSA2ux8cGRLclJ0Xc2OjEi97V
Cy1bmRNH1xH4l//rOUuhUBbB2jkIgto/bOfCuMbGwmUmjkfOSf7xakKjwkzCsAsz33oVSLCwnkEI
VMXSz9E2g6uyi9MB7Cp4dyhy6NUNWjGRNbGn34lmUUan30QGrDBEWLzy0T145rzTpNK0bdWc/dsQ
zS7Ej9jwW2oZ9547esBVhuU5oKQh08oxAmCLkIhxjOLMQmGtVmsRFlW29cx10NQHU4VCmw7ZoLni
Bb2VCnbyLj25RMEfcArc6UN9cs2DDaZ6ZAZ14QHtOs4BohXg+rneCMnVTmLmshvFF15T8f2Bc30A
AOqWsZm9vMaqFVM5+M96AaQGmAkv43w8AQ9/I23gSjNRAOWOxaCLLHQnhUDkTCb/Hl7wY4Vr3mgT
xLHELV9hMWTyYaoz0tBLj3jRnHbGpM9KoHpSfnrNWL1sEHfVc5Rc3PxXZETIbPyfja5UqWpNaSZi
OsbmIfqWGiEy5dXzeIkYmHEsOoYqmDzYelCrfrJjE/fBytA4XntQ7pSn8JC8fwA7kokGagk03bXg
PfvOJa3F4g032XZxOKThMhjKosWulMw2pBArd+eEfgFhLTg75lwRvhg+Vc4yJtYJF//lUeiUm1Ls
IHen9qKz4w3hnm1RsGF/UZ/9QICqJwBZgqbQh68MHPZ8LXpLQXBTTrB73U+1BZZ9vJoHM2Ek7/CA
BOSXwZZWZtEVewr5WsQ7zQ5+PNz1mqRpz6tu2KgfnkMta0QoLmxv6h0Lm3CNmkF0+QLfXE8stMnU
bKU2MKpFAnjK60wuDahACdb+DRp2wj6g98H9jxBqODQZjFOHGja2+1p1fJSD2HlTYEcRT84LV46c
POrDXL7xM1NRSgA+SwZfJp5hB4IUO4/yHtKDw1ja6Oe2Fn5yQvK8euA9K66qPT0NODAk8i2wRWmO
bui+byVHrJo/otQfHilom+JaN5shn2pwjAhnClYfA7Md4h5c2qXU3V78KsPN1ZnXxXfvQP4i7ykl
pKchSgIO+rsUv5rr8hyjdQKwnGVR4O5S7qbxN9eLrhVTqzCDemxD8+LIw+9KxeJRizib55OBtg3v
r6v/tQkXe0+pntO78B/38rjThwHKUUbOcazlkA25SrXj5LPL3nbIyn6OfI1NsyFQQmw37gMwh4la
Rn1oGoYwuEbHxHCViCKmhPTqOeJor8fKiMwXAJbjBtHHxD/3amgZwwV1/n5pa8zND+8YiEyLEJq6
yLM3LhK7MKcCE4hSIxiIdlVNr97SBoKxYchhpjXQNzzUGWvDuQB0KU26tRxACTgFOUShVX+c+hlC
2pLg0LZC6fUrq/FqqtrfzHPensQfGV2lKdD5yHzxni2eotnntzU6JApXWC4HIT++JdAPryX8F5Hc
cwRo3OBoROWhT+XuSqgK3M3yzVSFUEVOhf0/KBw6HUC8FiPIOPA5pCRci/SWIWc1tN2zrjF7BpfB
APW4C6t98QyeWCLtByUgzfV9p7IH7tgKd8vdzLBY5p82lCfNHVmp0slbj36i2uoJyYMQn442J3oR
l3UiBFgLj8GFZJbmHgyY2o44XXQSGL6CHXuh8d+twkcyBmJ65Sm/EPQWlW1nkUEwi/WMyIpUrYSu
MZExWzHf9CYdA0DBJrqsoe5w8ToSYbYzeLdiVSjid/QxFU11Vf5/WEwiIWK7DH/yqgTaoy8A/Pmr
rfDErbC86E/Df08cdGEmas+f9iS5TAZZd+qXLflvM0QoE5IQbam7M2sHj7dPigR01K7eFGmQias/
UhMD+k7fFU/bCuzEKPPhoWmQ26FGSL12nJRwT3pakhqLyaDWUrHLvkDzxJVa3tO4RWqiBIlY3epj
pCoEhdglnhm8lOP5/nw+RfaIr0rqozszRSSqECN15LAMbPsiB9pThI7gwWR7SzyRWGtyrZ9X24mB
Dmc0sTxshuJFKdw+rxqRAJbcWqRbrw8MC2CYM/p9nN5MGnFxi+jKW10mGikRPBPst1nQCmyM5vYU
CU/1Ly/+5jGbJJ4wywb6mT7xlk+MnABCitDgyqfsE+Xfn0sQpn2xDi3FBV3unkUNGH4hHGea1iSq
BlV+yXsbKZkTP00zTBoh5XGnvuh8L7ya5hY+G4AD57TFhJW79XJgrZYPsopxmiWYzRobXh8mMZGd
ps32qiP9vfOA56AusphRpyY2HwlMIXKvIEk6w2v2C1KGiDppF42xhul4Q148fG6+jvqRQgI19q/+
3DUsy2j7MPbjotmeRQMd1DcDN8BM+pnMK+2tkEuOEOicY0nNYs/LUnjhBvly/3tB60/D+e0qkUXM
eccwEIz63BM2YkiDY4psQkSV26O4F/diEkNjSbL5Xx2WDElrPOfgHFhxkd3grNPpGmU9x6SPFl14
ybN1YC62Gzb0ajdH/Zg5CZ5uW8cY+S28SUDLUgC8A2AWHG2GDsXQYnsTKKNxPP29iMPQRceC0EsK
ivp9+kEPBQhiT8r2bne/BodObv1TweTyJ2bRs2QnWIB5tLIR+m4YfDdhSKTCmAmXetf8Gw4Vt3vp
prr5gGmH5FPenO3TPc8eAujyQLuCHwxGGFHTW7wAbxttGv9bg2ANrMR98KP31LFtdfCXJ0ZdwHKS
bZwypzFKrxjQodaiMP7i0gpT/X5S5CSOCJ+wFYjYVu3XFY87+I8vIzYSviaJ4C0XiF2ScEqrhUBa
Wr5dc013Z8ceWJJlVLJz8a9BIcbFYCQn5SYuBiH8mDEaOz9JoUVJUrVfXbo2OI38O+K9i1/b0qAZ
kJSiYHpKFKPy4AT/ZDyN0lS1n/zsGK3LLZ8ldBBe/SBiqsjxd796KaImhoZDIAIKHp0h32wm1oNd
6OzzX/bIoF++mvX5QHdPedluPTVLTpvqYTrT2/kuHwDAvwSjP0G8UEEvdFeWhHwc0jbLSnP9Z7vL
341VQlnq9phrfaNL8YWNLrUceGA4Z+qVJ+W4lZPZ4BxuaiiszbX9zXEpc+0c5zkqSy2pJHqjStau
R4fMjOJsNCi8IWOketrq4g5wa5y5jHpiXX0KMWRLzgp8MiOe5XQUa9pAJjEsnFWIndXlSFY1T933
AIySqNJYA9Ra9LAGcnIBMlUETyq1KZEHuuCTzhUT+ftW4MfXkBw6FEGHx6dJ775VEUqvCHVmmwQ5
SSv1x9CsCWyn/5slSIHT/zn9ztG3k+krapHm0d53lPrkfxY6R9fiRsIswm3cKgrgzPRJDzATxqR7
Gzc1PUTC0S2ZtO0/7dV9F0Awh60aF3mmmxeRtNhbUyn+mwZosDP5rSZtUyu1xCX6IZuako6rtk4t
ogI9bla2luYev03AoAKQ+zpbM9R8nQksH70CZ9f0/VHj5PWK2R8CTML9XXJwj3HrChVfDtYiDY9B
KKVIXvu7JS5iCRMP+bDqSk3KFFO1NV/QTMvh6RNnNXC8e/TsBjtva8K3jiFet9XyBwohnmA5cKIK
sqIv3zRG7Z2mGS0livF1j54Gt+KUYr/vhk3jWG0H7jt3tTTBwtad/Ti62aqYAdv/1SG1DNzihXmz
bJXZpZU6SXMnL8tuurYSjAImURauroH80JtqnhnqQdpulhHJ6hIu+XNWiu8VRpYgsrgRyX+CcJC9
d2omyvVTFp8XdW71tYPHaAUvZFPX5owT9DZPazOUCp9WqKCWDVhoj+cSXNW/6XyWUfsNYM/hp9Cn
o9OTaHtKkiy3CP6SOaeXq6rTOFT9xPISI3DsyFvXp8sEi1v/Vx5s47JkPjEbvPhYZifJ+Oj8Hm83
wvkygvyxXLk7tcc/NTunuilAS8kb6bHTAT5XkdZrhcQq3CZYKZvwCuo7bVc5u5dUxlOj+uhOYZqs
sI0Et4ekPRXtCF+hgEcN/tD4MJV9vcuumQDoQN/c6UvFGYJozPOZDxcylRRIu6tQjocyoFhT/D1M
Od8c6L0QhorydjqSrO5Na4H7udvl2Tjuy1J4EPckp34KwTzT6hwtelxToV19rHw9kfZ/tqOqUpOT
/U+dBO1q/QZxrfmEuYwLjrPjBP5F8asPnL3eFmGGmdYcxcZoptRxydeYzczliQ5Z8nrF+oM53aml
53/ddZZJuNSeGW+xDSMWgyhemGMQh1Vrr7DFWdPfv9bovsUkemvuz9yNx6+5vgEDGZZ9+5YuVvWP
/VZaaJ/IfbkZLiohwTijwkDNru2MiCePc2rzVKoPAgBulqTM8TNdSMm4peWFFjusS1uy6qPkXFI0
XnSuwfQ09LZyfo5R1Aycmfo7jIklw2/GtJKitAGnKeS2Le157PC6rSe6KRJmqNBXt25A6p5arMNW
lMEmihdZ6sZgEb5bpMs+0CmpDDISnVr3UhtcaOnPhiDOeWo5gBtl3JZas2CelMAGBmkHIyB1iD70
UNOhsDgxZVm/zG/c3WvA9ghQqqMiaJXuvkutPahj1TqsUFke2p5pubDmSL/ZTYhfeYccWyvEhc6x
Pox9F/J2REG+PTQKgG31qsGEdeis34Xe6EctS8iLFqPnNs/KqPgdA8k2L6f8P2InkrSGnTzgoVkf
HGYfrJa9jjc7dhLCa6htElKFcgZBPQ9IN15YBjItcKz1MbGne7hIxq/E1hoyO8RJvsk09HzYa6VU
7pT8mCVeup7VRKvQ97MRJYLJLPC7XdLLj9McvCWYoGRtRff97mzIiMJZVQbNariTWqeUskcwLAKs
C2aEmLD9FFB13916BGZzpNdtKyQbiQt2Ywc5zXOWfGDSgGl+pSRm1Y5PF4wQZGFtn/cuw/DUw9Kw
MO7dOCgL4V7fd2ezgeTVvCu5fA5jd2k6z5svbS3Q1+pc+L6Q8UvvkU/7oznqZY5XQCLlS4zblPxq
oeMYKVTgkYB8WfAMZutbXGZmazliDux1aeftMOEZSopzhvoCNE+l9g/1hqBRpYam85rm0l1HwDrL
z+OSACY8WVC/NSxxwuTeVWfYVXtkhBUxOKXSqYQKf1BvonxpOe/pZr3bLmGKxgjGIvgM6IDtV8ah
+LW5ZVLyPeuqtHnhSTFWTJp6TdbPuew9fkoJHCyAji8GbgfAkI6EhCjrm3B269Zm0Xo5iC708ady
YssgAPwBJtA2xijczFjVYqUqqd8CRdVc4EDHE3iCdjKtWieZb8NUFuDrQcL6fnW8tyo5fxTR5/yH
2eSfjx8ieLOHTaKW2vqm3sUqZ4GWys09xLbvMwYyg9JMGOYtIZKxbff7Tnoc4omwmRsu8f9g9lq+
M9m/vm037wHi0YZYaznl84tJW28DNz15oP/DHvYcprLM9je6/ygMSW+yd63x014CKVctYOIbLX9j
p6PreABNMp3VSdnVw5AhERY0L6gDNZMZ/XrUw7zaTf1ScyW0my2IZ4rUz8BsBEFVQwyzise6c9ra
Y2heWibmlaqqN7LU+1+/7CaMuCGYBrsitMmNfGQ4uMZVzmBhxbBflvklJNzJHqyZw3NlwnwCDKZG
pNwliMdBQgkqBukIThzUlnOx8hHtY3w0De51KV56yNaXwR8Y23igvZHL8lwCkiH59tzRcV84KRTu
/fUChPKh/CrpoXRoXG3R43ariJ5AnGwdNR+7TJ8xiVv1/HuuNCCJoHhU/tJFlYSmdnOHUoFdp1RL
8NBEoy/dyfZVAelfyb4wjewvCCiMp8mJfXL28sZCd4t+xF5h6Rz32ymsOt+ZMwF/wqZrA/QFxDay
nDjLZ5r+3So1uQNgkI+VrHcQS7qS+iekRwN8wJVYrLuvll96yd5kDWv2uLyiqqwJEm11TFb4x2Vu
Fm/WqLHFoA47OLXTnh1IwmQn1lzYPN+lnRIv/Ns7b0osaB7NcEoDA7Tnm3Nn4zwpS7dsckZvFGwj
rmpixtL95qpVS7chgrKcJAfy6Bxf6VLErrIo9DiQtxO62+Xlo5Lm1W10y8kbP1khV+N3mEc+oY4g
/eN8cY8nY0rz/YDtpcVVvJSFY237Ulxr6aiKJD/4GVUx5+kfOp5Jxtz7FdvHk1D6aUS8d2Swq289
lfvni4oFEO9Q4i6d9h0IR4+3T3JaKa05+D5sG4iHXSr/CCnxCe8Ylp1RgZEQFPun/JHSOds2vjh2
pfj68+QxBGYPld+qR4DAJSKVfSMmdjvMqV5fX2XUYaZgXsgiRQHA38d2rXwwCiKnndlf8O9nScq8
o0hU/tJhJ9UzXl/MdElCfiQ+HAsT0znAhisA6lgjrsokyv0FfOPp/IpHNrn2/PXmfSYstHziFj5w
YDsX2adnGEZ+2kddQqJq0qyCML4KdUvxfb6GrZyOmkZjFM/F2mHl5G+yTmTcqlrtL1ZSxpYD9yPu
DI9WBBHFYdv/a0H0oHDJdmPqQzOy3eZYC6FaG9dEAgPbC79oU9JgTDExLrRI0PYwE8w7zcUWZ4k6
aIjQwCJgG20UjbcZNeJMSsmw0zqtM1ER3rxNXd0oyEs/LkkZisGVcNlJxRjePn3OuKj7I2c/90AA
RSB+Igij4/10yKG11BalAZUZiRYozS3cxpLlzw0oMiBTlacGB15BWWh+wzfFwgwCF1AKoqJQT+z/
Tm6rZwo0ldzVOWbL9BkGhxHDrqRLU4jJTEHBc7koeokJ80PzD6/sYKK3I/TmLE64tANovOTCgBWx
TZ9LEGW76fI3HUVAkum19HvZhlBbg+UTypPOEGZDZSTC4WfzZL70gLwB78LdR+KLm0SFdUSRh9a6
IzGTUT4FTU0CWg6D5ADrfCGK1/4ymQf4RSSZ8pLXeL+X1rNQO9Zrtnq+iZNsYXJe+X0hZJGMM3dZ
AkI6Jeb0RqSRjrmctnih2rdzd48pX7MBUKJfomt1QijdAECepwaNwuL1RhsM9e/42Si+SF3+JMrr
Vax38wjj4nLbV8OUHiqLxqZL36rsCzPmaiMhrW+3bPQ7b6pXVNOGFe8BUXlnGGUMQHr5wgDBCGMA
IQgF1I74506NufGmW/qTXS3behQIc1EO0C5qkYYuMdWfw/7tVK7U38jqM8Zo4pjGzl79FQLlGpR7
TmyuUvfTqZL/HtKy5vsdo8TRCivuOBscVuAYkxHEKiUTNsy1EO3w/lUhWNkeBO8orY3opdPOvlWz
eWyzRDA9T0LI8kJabzYhpkc83TO/5vXeQHGRtlu7Yz1OIuyrrscb8PmxgYk9uX4Pn/7TN+RWcogS
tu1Tir9dC6zJfBBM67nCQ+6wqTht5O5np/jSg20nzHBVkeAnCuMCQ6aVZI9tJhRz95lKqx4fA1RD
0ipypSHHUeRb5Zml0IvlptMmKvzp9JPpD6rqYuk66VHRtoK+OtG2YYlom81GbL6SfzJnoXalkgY8
dIv82fsX1vppYxrEsG1zKRTVR7kmBxLDOPV5UBKPhyJjR+9vxTZevr13mI1Bo9Nq4g6wc1POzu6X
yY9K1Gs4U0+2/e8Vd8XavlMsJqkvKIgb7mfMn5bJbacNNjLO4zDvMvaoE/jC1Bo8YFOJQzz8aWS8
joPFKAQub2yfzw1VkyeYTmxwUYXvYBUtPt9n+BOG+8AOS9pQyN7GdAVHCGAM6t1eTA01+WagYo9i
HUC87vY/Acl99unULb+FUjTntvMCP3t+aXYoybW2W5HdOd+AXjyP9eyhT9jWVtRtvaJL58r1chB7
zcjecEpUn1V5O4cp69aqTrDYMkBFXZk+rRzSMiHtYYmwP/9JB5kc+/b0Irh7goZGkrgZvJzpTMPk
+F+wbapGdx1PFo9NXQLCfmkSoF/4yfMI4iZCow/JLTzrVUQj+45LqvQtxgiT50we8rdqmPDabOBt
PA6ia+jMaA7Fq9bb7KXLgwkLRW0UbR4Y3uaWBtKJRbyY1wtvJ7ut8/Uai0EFNYDipz4ZLBjhGqJT
q/V6l44aunXcOG8khafaHGjD/CnHUuMakzyGETdb1S95IHb6mAzH486FoknU5AqDXGcRASs0m/nS
pGrBz/bBuvIFc413aRpr7+qq91crhI6DLaNy3o27lVpRnhhOgVCNnBnI5flezQo1/zfExNfssWQ2
RPFAt4POfmsK51Xk6KB5KDjfKRu7hAT9L2Y2TrmTogVrITHB0Tw4Igkptjw5JOQNHQHL4GWh/SuC
xKzL/sdyYJGPI2MqhP0fexeoC07MY9Tln9GdCUKxrf5+soT+21M/yA43QQL9v1C1RM01/1tMqF0l
7N6PjqWmQt23v6d/oL/6NHWgkjzZqaIXD4noJcrbYsI2GMlZe+IRRnTiEzrN8m1jhGXFe5s5trYa
oexcnH1L1nSZVrkQyG/dfV5RUqaxPFtuVndKhioOpju0JTkioiwXjKVdCgyai0Mrkg16yS8RDfcj
0Nw5wegvhAiM7sY2t6F3U3/MGG6bwe0rrxE4amSXiBtxXZ3V6QUSnHNSDl0SxIZpzf/ZMPcpWhZx
SeIZ+T7/sM5eDP3nM9oGi3Zf0+rCwpjJiK+0gCOMhAasz+sHhItKEy94hcthUqsWjb8Wp7pDc6uz
gc0NYRTSi5tGpGzcGPnNIPDyvG/OblCJaz2UwqHHKzSu0D1QuvuHweyqiGBL1besDfPoUkXkURve
MQMkYp8A0qUkjcZxnaZZEL00NTpSZO8wjKLhThzjj9lqyIt2iJqEne78yZ4pM6PkpdjYSvcqL2b6
ShZUfIEypTbQO01qwyz6/FWZZBOHNonHoLaqPKmu45YXeLjgfFVUXagGjtUYjXNY1TtYk0QQNw//
qHlI92nn3z89Ps30VocGHK2RrRyedkyiqsEYQIAJVrMuxuA6cUu2gAF9QJf0x9y8yuTx0jZ0l4Wj
bSz2/gJGKh/S4qUt8xFGPn8GNnKpbLoTLWnjVXZOQ9lz43Pr8Te7daAJaEUQZJpY8RzAvhcnpK5/
CVa9PkbdRDLP4r5G5LAT+oD8B5Kp6/AL8TcXI2y8YvNbRewKumiVCK/l3BjA9VwKVvBDivre/m50
ElSx823r1HINEU4a0MbHxtzy2L77E9Mc4sk/9YWIZRBD+My2lfsL99B1AYKl6N1FvIyLQ8n8jo1r
mh5s82Gy5Gqlaq84+k0G+8KGtTICotjRYZniUGtDym7xaQjqjheTqLVSt5R2OaNggZ7RDVfRUhty
LHDDR0737obPVbrFSflj3HTk3W85LIsLnD6Z2Og/fmUhcOgGrKIzOpik6M618Dx6CoTGPRJOoEnH
xLR/OQMv9MeIEy+1Brc+/TOEY+2v78UKAlfoY8mfbLPWRANVFm6auE5HvbdUcWX9tNQhc3iKEWjc
Zf+Va//sPHZIY+/ib/zvEZAN8bFyOjX1gsyM7t1qA6UF81XfNvwp+4amv75S5RTbGdBObTuKZm4a
xeYYON9RDK6mhgl+cXhtX3JRkD9iHHeiz0+Z12Ougze0ST8/wHTABYsf4ZTwtbLIegw46vD6M51p
FMQCYNFK6uGy1U/9ra+sltMRZ7TRfCbtkRjfC4iCPIRP1PcK62Wg57ZDs3BDzdMDAFS4yKSpltWw
hRPfkTXwm0j4k0BDTPj58/JO2xNxMP3I81/6psC+cnA1tawIyWC/4CpVzILQpdHnw/wB2JgRPjAY
mjJcB07L7/jjy3EwOCO9uDxLcsJgTnSbhny7/jvhSITayqhUkdEqL+5H//KJvCL+8vpTx5km3o6Y
ZkfF3KI3viAUMpRhh1tWaip3M4VR+6KHNqf7Igiyz6X+2F1pIm7kdwdEzox8Myrrmj2MXABOjdqu
Hcjs+zg0joZo5zlfYwFG/7Es1RY9cwbEXjT0nJigzUmedJxEVQf3l0PLBYeUzHDni5V5ZjzcRrFJ
E8ECBheBiGcGW4JaYXsiustzB6zKQEtbT2OIZmim5eF7AtQkWxBShstV2cFjbMcJNOHHdWIQ07xb
qkNuYr2ft6ayXU8ZmA15+1K9x+PvFkwXV6B9T868ht3ZgfgGcrcRFkz9V2abx8pCrOf5FkAal0Eq
QcvyDkiTify9BOEcdI6/Elb/jBNqEY12/5lo+KqT0CBFo4DfjmTHWUix8hwv7ORqZymqzgZleGq7
F5DAItMTXESvZ9iMLRT8jg5xW+sNFnds9Rk5LiL6xyA5e8Ge00zVbVKKCzDqLjleUA1QXVQC8Tyk
9JNWV32rBkHIFdSWEQwkQIzXgenz5ZSBRBlJfa3NQSB/aE6rwYNYIih5YkfGfUNFPJkRPCNTEZPF
d1dBxshzziOgxzCOzMfW7vlONv/ZuG6/gKZtRqNmZd1nvhrPSjeOYRLV0l4VAh8EoNGZPOmy9Xxu
1W7Xg4xDx6a83LXKD0Khj27ZmRPpZ7rL4KPNrx8dSqu8tUl7VmM1l5QzU5rd7VxPPcjLjn7jZXJ8
+g2DKI/LAvKL7tKqxs1WHO2lQC+FOZCLDtoloYV236VhObtMOmFhXuqmW8ghAb0WcdLbvsH41Tmj
yiXBjwkNVsRPWe8AkOf7QL68pk+OWgN5o36PiCx/ltfZTtvrzGcNRRNF4Mbb/RP5xy1IFMBvK+bz
fhYu2IPlqWl4Eg4K+/stupmjF/UKccqUVyFgIMs6Da6IrwqmeP3FYksjqvSvscpho8i2qjZWWWM2
vKqrpcAaySyyRyQtfo9n2IO3wLSeUgk+xQSVvhXBrFgnP0XzWU/dEfu913ehXl7ENX4pzO3RTVa+
l96wTDgbfCOwZ9DwjEfJ25JeoIihnC1Bd4hh0+99/zJZ6FNkjG6SulSiMjOHSGyVt4oscW98GmLS
B5CIck00WJonZN8Kn/DnVKCWAwU5WKuzCnYldCfId9MibzPfXSolngZFT388c/q60tu8pVzd0kXb
h0dS6hsdKjA9RdDtpbvAT3xqhZ44RhFEWjK4UGguTC33jwr7vhNIQ6DQmah13LsLcnKZbwaa16GP
mGB2dGjrR+pFGJkyXpihS7nNGOYPPmdXYq38aAFJQMGcexprrRNDY561LDJ3SsnSFz8RVA/LFfCp
r8Gd6OnPHjo8CrORjRc7J4hZbK8/e0V7kFE89iaPLF3qzhYg9RKmwWsJ8m4I2rBozJ/A3LYjiaby
9DFPCY0+uNBnoZJAMzmllQ2ktQRucUygSCA6plgGJqxuHgBAg/1aeZq2dMyXdtXnbSolXn2+ioM/
MMxsVuq7pnn+4E6dvn1Hj3t3P3yiOGxzUBGIosQ2LRVq1hf/ZcEy6rupgyRap+to4fTAc0rLq3hx
JEjavXsPkx3bv2c5aiz9t7CT2LVidTlYg+nS8QG+H205NHR9DDwpqMHvq2b4W0qTRMoOTpjYVYhT
UE5F526iuEPvL2Oo2N2Bbp7Hp+MsXF9Jg5+6pJ0UQjKMyPbslslU9M8Jxxo/3oMrCIVuBp9i/pww
43XF/zJxGoMqByS8T9niRG5ZdtH0J7of6grT2eiOxkVTT/opQ40+0ZCUctrQUKv17JZcBuV+VnP4
OTaip8ucDNTvKmzpCnyZd5OhrHaZRpt4iQr2nbXmePfAZKHCMZHJfXi1FTcp92/Tv5J+BihItp9Y
tdSwBnLEcCxoKGUzA4XWJLL/QPrUhTZhWlS0vfbBsOokp7NTZcMiPGsD2Qz25mlXby3oPFyBd+Oi
zNksWu0eYr3nUBYYOQloquItj9Pyp5O++OPi/b5uxjHtJHhYbanTNlKNv6UFrIL/hxDhieMoA1C+
9FQDIhNL3U04WYNiASZFpKmZOXVR3pmgFf9c7Kl+fUL5LrqA/+GjvlemBe0rUq76ZaFn9eDqKPIS
z7ECbbrw/XPtJ5kaqWpZFMVrCvjAK7Xg/yUCZZZe3TIS7t89e+JcV73/fyFricnzYHYSjruh8Wqh
3O2f3lN8TGXtWmSVvPYKoWzjw/mUG3521A848qybsnbA7tWpCezfrbKw/7FqOyeK4j7v0NDnbVCY
9RDqrRHoem7dRw6ZTJnTfc1cXuvg3SsccEsHveb1ajsZBulYqqTKFlmFFMfbiJ5KO0zJouwAcZXd
BIIymoBHSUeWthKc5Eud6Y0V8J4aBrmpkCZaFlcW59wAEl5ZWnOeaOTAd6nqdrx1igOmd2BFHFuw
RYX8gE23Tpsk0bKcfXvR5Dy1JxSYVxF9RGms3MnXnjjQuyufaltN3fV79Izx/AVSlhuAl7zu0vLP
0JPepzaax5JlEkukSw0/o/DDn0omS/Y98XBnHJ4FoZY7YXK8Oq/mwXcGiU5UjJalyt1avQbafB+8
kH+e9jKFN+40vfUGNxy+upV4bZPN2ZpVrHkXsk1y40LVqdw18ARzmT1MeP3wszfjOMuKUqMjBhaU
4OhChuFM859nui+FyKC+TOCuJebma6bNBgiCdaPxkg7hK5P7fgKdaJyHz9NTu2YJxp4ngrrgaNXK
vOp+nS8MbtByGljhGQx0/MT+6ew3zkI+FMCRLNafLkDhHW2p1ReJ+WmAAspn4jOxb1bS+COjUZFh
gxvnpeZfUVjWhd7lartj+5aUpv2o9auN3lgpGK2ufLWK/qznHVzir4PAmv+lTA97CO1rFNJVpmI4
M4dSA8qbO3kxWaVf4ByDtMKTiXJZMLpYivW7MpPy1/lJBjB3HlkJaan9i1/xU4ji2tbuucRuWZHN
M590TqqgJZexy0n8vXgsGpY3MoFIh6bjGSZklM4q+VfM9IliV0HDo2zGpDvmp3tXYUMsH2BowdJo
ejJox78YTOn4ji6CmlJm7b3hcs/c/x8ymnv38Za/aIb52uw8RPMJBFrRPIb94bgd0pBtWS3RqWZU
vMkY3B8AyDNDYOmp/HIEo9ZTXdQ0dfEtgPllMtqOpqJ4lCyz4SKSyK7bGeLK8663ZWp7OUmn/GEQ
eU1GUkIaSLVa6YUlhi8d4MEC35MO+MtRRuepf8bq1B7qPltLh8dDG0RkrPP2d4DByOs/jqjCnqth
IhslFVPO4TeMbzekwSbcaJ+wLaQk0y58PN5N4h5nMvRFh3HE3HNvi6UwUVQBW4RjoAqtrkWeubUS
crFSclmmZ5NaYXxArAAn7dX8W2sG7XH/KR6Bgik57CJehuIw8Pq99YqDP5fjzzZQOmOau8xXxi5T
sMOKpWR2DO0re0LEOZmpLvhmUoxchrGqiPkjRzLVjOaD3UPd6VG2vA8XVRG1oiwkwEZXlV6CgADP
9faI2knLIx6zD82DNvujb0c2sHX4/qqAzqz6HvlF/5NSpE7bIb7yILjWscJ/mYyquoOOIdgymGRf
EBXMSpQ9V1geTP+E5tDte9Ls4p+Ax3RApmz+uPXs0jz2EISvmSrw+hZSE1ES/g9WKgtOdH57+LbW
iB+GdjbBOSD5fwzDfkIxQMhuKSoEffVABbwZ9POUmPQfPmamFZTmLmdkGN71IYYZX++H1+AOClUn
CwZ9GkhKlWaviN6Za0DgIjZodAXJu/ODWkE1zsl9lfQn1dlF8wOcQpaBAB1suRFYYBt6NqPj0tA3
IFYAgM8/UygiB5SHrY9JmQ4+bk2gaKS7Mhj4X4H4W2IJZw8ZZ8N71VXryzBI3n+oCy1jnCEVhn85
5n10J1JFCFiRdNqXrGeY+JD9IcH2DVqFHRLg2NEWnR9zFaIjZ/meCLcyZ7Q/CezVbrNHBrGMvOYJ
MsiJ0KuCD5EHTm6B4g5GGInfj+mQ4uKcYl8mk5slRgDGBAJSu2MKgTw6efI1dqrCXKSab/OBo3Qx
CUR3ORE93yzYBsJBQsGNPLbHQo5CT38KvJ5sWM+wtTM+JjOI2fN1wniEoYSBZv1d+MCwYVhLaIK2
EpOnPHT9hVFD9aTxdAkroMwa35t5xGi92Xmf2GCVyktT0SKjHlD2GeXX+bP4ImrYxLRDPiCZlBJ9
3o4Lakg3uJstJIIEagOhyVm41PAh8wSKhF/ZeJCy5SH2NLyGxST0FpEjC6gkb2BELJOZnHfU63Em
ZgZNLhUHFpHYZMxzlp4NUf6O22aA03l+Gnnk96iUw752BZ4ArKk6ZZQkaW0ocgc3Sqs7DUEiP8ZH
vrxaASMqJ5pOZ9nCpC+57twBXKarcKPprQKO8AfAxbpTtA8EUB07+ulWoELLJMzPo04luCj5qI3B
r+20HF2uceuZCVe2zPwlL43EcvGvUu4vKV4BxjoVdaxlLGTKoWxu7rNzYSd7UyaaLkpQNb4X9eL4
du0ANEu+N4MYNMk+MnDr+DyDbkMaOpbngh8gj13hdyNS4KkKSwpP9+8mbMpl99qbYW/oc79cJwPh
4I1qi9FjZKdwC7Qs4Vho5NlLLQbt/HONTSnkVDDltnSmttJOIYoadVs65Dq+YO28zRv3i+02YzAg
dcEaRr2Cj9RdP3GJ03zsVozfviGBkrwyqHdBKdi0Gv+QPygERjkwcFmgv84WJv2lJ2GzhqzvZX0P
56a2PhcPSfZTSoxfEz/hppItwABmiDIds4B/nG1+prWpVOAZriKySwd3AIRcgTVmLaFtNYOT/Jsm
JXbc/zlKlc6mOHrF5Ntl7vl1YUIZ1yvJiPZmhqrKTlL0crlH66TG4vsVTkfg76KPNRv6nrw74B51
h9PztzHmgeqgLvfeQWFx3V10McVpOyPMckDR+a/jFNCOx9YW3ahaoQdYtV08W9TWU5VMhRfRfvkS
OM4Or8hSRs9oGVMDTth85F77lWb3O2jamQB1h1wdAeJzz3QjooOmvZvBJJwzbsIwh1bE/GaTb0/l
9qcDqqws4GhguBh48BZGY2NNIJeSfxsz70YG1MeqfKT1muL4/9pFr0+Hbd31g5HVGe15UDgr0MZD
pTooBgP+3oakv5OlDFOJGf2XwAxivvBQ6mf8bxxF5gTUSfnXQzKxaz4xbnbiRpQY3ljPDTXxCSws
tKzRmpZ/SudkacYq1Qrl7hTt8KGM5UhYvoTjF84m6LdJUouEYTBGE0TrBSCYaugLGQj4GR8Smegf
5fVBAFe1cBOr9xYJBB5C2psLskN0Xd0MvUf6F/oCToAqgsi9+vH2h+KMUJt1ORErLIldxfGSYDJd
2eUuDUUQN8i+e8aojS7H36DiA13Xw4L86lTV7a3UqpvP7v7+Sns/1rWL3aseRsZaop1FQBvMuvt4
fAAYafw8hSULg3ayq2d6o/g/dVqKr2dAl7ArJBTVbl40fZIaN6SBQd6FQGLISSAVkSREa1+OXcmI
s/2nqal92UP3rSfPEPIlV8EWA6v//uJGvhnjop9or3UtzkvMlUCxjyDytL/HUMezdVKwZbzbaLgg
LSwZfcaKHFY63UBGGqgJnlkcLiPTz93wvgbq8JnkP13XQnb6c3k4XFJ1Zqd+7mY3Fwn7o8PRSt+3
OwFdIGCcM423ABU5yuzrulBGZRVV4PowZ7/DCPuxTM3DwihqzNLbQxQlUDp+TzEscOqe0fsYoce/
LjmBE31V8dHp55nZZ1ivwTOrmOC0hldf2wh7XfptIf28PQIUecsPGlcLqybp842XWUjKHUIiHwCn
3uvwvUR8jQBYI1rU6Ux1Kg1dENTCSJ0cY7Nmsvb27PDcdnkywWVM9SO3K2pLhCZV0zVvf549d6b1
aZFv1j9ceq/78T3qqrvp5rxc53UhLngi6kvvIHAPBYyKhppv43DXklh9AM/akDeoxdyGKUJK3jPi
gRKDxJkU8/FIQL2jAvUc5xcvgT8amWMZ1anN0RMKAwcsgTWchkgaALjZjjSOCsu3lq2zqgMzLH/g
EFFrckiR0m0BehtAuOtoWD4qCF0+XzLouONROeXVTEnt/B7Kyz9mR3GNB1FdtJjNF9FnDrxZvCti
/BJiJGceJsN3S/PceEIaaIsgS2LtL597pRc2HNj73BmVL2ig8CeHFJnpOtoDYhiEGpSb3++D3uBD
PtAjzWNbE+s24GfYcC0PzAj8fhdDGwHfDxIZjOmxnau1mKgDkDhu/ocudsletMjP7L4sXYcD0mai
x2ezIjRbQQusQlLc2wI4tEK3fFfM19Eh0+An7K0Wvd660mfFNDL9EQdbsveA5rZ1itciZHSLWbsb
MFZD1YkAc2TiiUtaGuCpoGdwIWcDXn9/9o5uSQ4E6FfAvbiN1+yirpGzSK/OzAkpP+DryeYmNEPZ
0HX/uHNQAB8Oqg7SiZgwFz3UWZwvdYn162s/M2xBRrUHx3WYMG6RbcxIfWlE1Pi/+BwnDUOPqWDP
EHYArtK6/IBnnczk9pbJIXNjszfEGmw7HDLOJP+0igs5lQCVHZsE+athbz4025ORlVceKb0ZAKg+
X6DTCqIe0RDFiX1lp9TLqGidE8FDAazC5pWjxv2EnhIjO17PzPdJBrDASQMQ5NsiAIyoThVey99X
wa8zpwk6T258NDbEzy+cc3TtMNHnoUrcT4GNoYSHtsyGZbl44Ta7ECDiQkpktPCzg2BpvSgBFdQp
JzH2elmCH1gYlFk5wZmJ+nucXXm+QhYYm/L3/Hb3y9bxHXugW74BJOcdPmOUrqFG9qspyYU4nr6P
qqzqh4/kSUoK1qmDtEeBiSRbNvu8j07Pb9TV3XW2ikLr+EGc4rSylS1pvxVEnbknPCoWx6kteG+r
kSWrN94vYYHz6lQsZUGFeZZXLs6sdpiec39j34+NIsfEEhEHptXeZxci9jqOumWVRNTwkMlqXBjt
KVSxqc6PELPY3YmjHiqJ5nWcnNbkH7bdqDsyOig8Hf7u4xbnM8C0GWIExXu/iJq7EIcV4Dig/wOv
YGlY+3Dni2adnQA38qxsY6pi1fDYnVGDzH++b161ORTB0geRA9Ouha8oKEWmR+fmxyfNPHrmcJxL
55vi0trYBRdMwGTn98ZOtf1/nFhYJ4/kZp+TM0G/CyuGRZXhiIVCEQXkVU6Mt7KPvicL254T0sy+
MGr5Q4mtQigav4zu5LDJT/9zpeCQjz6mKSB+Zs4mELmYFIfEYLKDVl2BQeUcEbaDBXlVtQgCtvDG
lTSjbmbS/Our/NI58CW4iyErP6pMQhq9VifBrb50Fq6k6M9Jq+3f5OevxI8/9Mr0/Dn8pX1PtKAO
GV5ma8zYvOqRSIgmHRn/wrl5fEKUEHW5D1rwpuRJo640HIoDp8GMf1sxWycpHx8Z+f0GjSAviM93
+JUuYO3VF0qdJYJIQQyhHFWZWxp/tB3Vsn5IgZygPrtqIBK3n383kB2UdtNol8xi3gYE9xx+e0Ew
FVBO6AeGn3/zKyoVsYZtAUdjnL+vxzwCUNB7BDkMoAN4orGIPvH4uRfBhTr5wBLk/5SM5gWi1SeQ
saXSGXHlD7diWLJA6GgJ/UA2eAgep+MXDkgmCZXLi6vd3phSJxJw8bd6I5bXYK1I1u7fpfbit7cg
RSOZSzqwms9I7pZ5EoD/uODUtL23sEalIVpVUg+aLDHOnSE5xuTT3x3rGUNcE3GoStlX5fK/TuqS
TMp2WcWsZHTQSwdQ+WGWISOR58DUNSiBPVR+w3ufxFTCT1JE4Yzhv/nBRObTmuVNqwQ6uF14178r
K1imcHJQjX2IGKeFA8b+4BG40Hmxn7RBbPpbrRFnjDHDihNfMe8qwbh8gHQKNuqp11+YNQwy41kF
/Ak+z1PEXNeUKhDDuo31jcF6ipC9Pk1uoY+ylL7BVfI+E5q7J0zq2y+AE7PrOW01xDYOOMqzGypu
OeCdvC4VtLQL0jo84uexSRwsHMH1qx6mOt1CNfElPtsUcRH/0dUGibNQouTd/SA2Stbh/gRC3Bny
nYBITe5d7M99OwZbr/KaORFu2nxeAN1f8YXspYZR96XOPY/cMKdcSRYqOY0pppwohHdaGlJIAHBr
dkM0PaXfOtQhH9Pt4KxZECsDtpphCp80a04o60Cx2+zW2Y3JzhUIZtg318ADBP6P+94EG8nHCJw7
Xb6cCZU6cXWaUz/FuRQnCau3iRQNDaX+P7abQQZM/1RpcBy8k280dKlagEp6/cq7Q4f9Djl5I2zW
WYxXdjLG22RLoj9mkG3kkxjcsnXDPu+YO8HqyJKKcu0UXNyKVp7V2pq13vGKHwWG8KirSZsLpZcU
s9fG0cqQyGPIixg+THahfWNuSMheLrHMLfBePE46JXqax9cZVdMQ/L5HrNjfDZn/rPUG/kM86jKy
4TI6F8bwJLQf34cy08HnNQQrsjXSWape1Z5+15XbB1v6PHuXCkDIUrT7mbLns7TRc8LleaZXS+M1
O8krLr1YFU7tOmceg4bddqG0R/QoLW3eDq3QBmwesp8eSgpymxx0lV8QpPU5hX5tyLw6+f+rbfrq
AMtl4tOmCv6LF3IWJlnYLvo+PBdkjInVH+jSkPcG70ZUhUa+Zip2oVjp34VPIDWsorNbSK7hPbST
4ORn6gK0bcCcTjTQ7WoGVHVcdM7sLCZQ33IcL5t3YuQ2kHvDbjWYdBW/A4us5VPDT/2o4a25w9Gq
YLSg/Fnr2fCqp1avVrCdJ7N2FkfAzerYeJYLb+kKc86oLtIPh4TLxnzwyY68fnMMVI+QxMT4ils0
EvOgeBI05zYLwhRZNXLs7Bokv5S5PCrxIC7JqmkpifVCNgIOt91+oHlGFDF0pn4bb5rJSWQxpym/
GD1AmZ76J8jiDb4lstjpxQFE2GF7IbqGrXvGxctbaf1PCPaNR0/2izRENCRmn4Ma4Vl6jQU/jbg8
U8Dm6M8zp7Y8bNehQ3E6pQY7eMeMP+fy7eYPZvvyPNOheVD5f8ywIDf7J0h4IDYg6IS81xScZytC
1G8UtDKVKyDf1wm+99WDMa7DtfzGykXBws129wnhXG89gY+ucCPNjdczjAnO8HWpD28CgIsarRyv
bWffsK+QhiljdG2mui5gho2aGlFMiFl8Ddp/ScNo0uosWIVsUF9Ffc5gG0pNNfoM72a2kXgBLn0W
gn98M4AVtIfxCIE4enKtGxB/vzfO/mXloI72so+I7eaIgAnDGgo52JYit0kQ/CQ1nAoBv3FcxGJE
/8H2ZgFGmDcIlSwswgHMmoas4pGZMz49bgLwUr/BzGIB64hvANju3SZWlBNm4zG4BomA/RAdT7OM
6ym23P7YXEWzlKct05YaHmAcNRLuJmXFZFLkcCQ1ruQwfZJActc5lvN/dDORsJt/E8bcsVlQGyW1
daD6MzOKslTPXPPUQECgdYmdkU3p6ZYXAxUo775Fr75EyA7Yw075ZHiraqLEEifmrWTwrz3XVgIe
BPk8dwAyYuim9f5IVDQKNVWNaNKBK2z2Dt66e+/CPpVGzbXOuOnOEpDCJhdsjhpLZzL4i6AJBJvF
qEEGT72yVrfJZ+o9YRsRPaBmjyAfELpvkN/FHwGMd4ZAuS4wZZDB8gvuSSwcdQNfQMWv1wJ4/Ost
zTX8NQ+XMzmhpLrq0V7NSx5ULBN1nVmd0H3so7nND0hdmw3ilVzsyLn4WZANWF3MQkUkGMRJ7YHp
sdPnT6DuZ1Fo6gEeoJUrr7GNy77P2I6L9T9uk3zYNiU5cyVUSnlXN68PCLcj73crYS7/KiwV33+0
6gMudBXtV6see4lfvlQCQ297gN3HwXrwv6wQYdG6ZAJKOoXJ53QzlO/myzzIDUhRHdi4AJCZz4UF
6PPVb3CHx7+rFRZt7nrKssEosIpD78uxLDrpoC5ZiJ4WhhUOe1GiQ7CNYPryL3c276rFvEAarQch
YvSucjSw1GSvHwSFQ9a/cK/mVp9/kxddV3OBbez3lHxTWKbjjgNmczw7Fv37Q7Jd4crO0lDP2tSh
QOeAM23cUuFLnm80kgWjzwyyvtCGPwuegfQsADRDNUJxMbDdTKiLFvgMvh9e9Q0bRz3/pUBy43Uy
vloLj5Lm5n3cgmPHCWflIBWnf1eO2QQfsU+IeMilPlD3UrH0iTbI98pffyor0Mjfj/8hOS/F663+
NpVXYcygnGnn3/GyFK6cszj0rtkEv6WeFsQWGoOfvqxaybvS47krTc6nepwUUx6XvezLV9dp4fr/
ApH0VOFtZJYDLvk40sH8LfkLz410lvAvA2QNq4y318GNg/fxb8M/AXsSZEYNdYQOEElHBVv2IHCm
2M2sKlRLXjiGBXPq3OCYJh095sKrXT5M/eBzhCO8Dh2ty2uI3Pl9rTyP/7sQ6gnuXv/8xCMuKt4n
haxCirqQjYjn3DnmH2IU/AQNcOyepq5aZ/wJ50vtrWItXRqcaWA6vUOT6JiJMyq29KPIrRXBCi2I
4r0UJTDRUIBSOAU7OkgaEaBsfcJlz9enREiwYamDBD6e9mKsO0A7BvH5/bT4C+cwP9lKLUalS3vX
wMggvefhFKht6oX3qwQzZOfWJQVZwSzUAdiG4Ug08PgS2+E9aLlOqd+mpKfqhv4tjJ9bcEzwtd/V
lbAXiB6kdgDgYOtuTzM5c6nypGrqQ8HAkCLZsUZc9RS+gEu1CmrPzTP6puHezdPXfzc8Be30Tini
22A3jpqwiYQKItPA1CU4wmvxe+wZd417NM3alz8GrxOBKViawSKUVDrYTEPvPSRVALkXK5d+1NJy
JmU8kY9d3Dmh/XOeJZKXhHIlxxWhqo4hn4yDYFLo85th2KvOcJcqxpoNdFFuZjcIAiOCxD6bqieh
rSyoKkTkQ/e+3HnpouyzJa5use9F0YAc2PmW32AKlVVtMD2tgmek5r1H0u6lwhuR834bebKk++eU
5PpC7srhdrPJsTwhKPSbs7d3rEEiLCBy6++kC1B79p8sCyY/h/v74OJGCVtygBx0Yg0gFd3xI5H9
Lo3wM0nBOXqcYlHHQ1tGVNqCrj15Qq3PRaEdwr1ukAQWSjoLMatdO2TA1PAmQsf/HMiVGrlv70/N
1mb20bzXvfIW4StLv6RUq9b/kZH2chEnJUghWJ/qM72bAtfXhwAlM8+dHaxzJfgnaUu9YTCJZzvb
ek+JWuRsnKkGfX3r+7bYCEyCWkoX6NYJzP7cdcU31YurqzFlCKgS6Lugcl5YuOo3irj3b2XYiJ71
WgpBoEi6cBg6rzT/7KsGFOvrtPVFS97R1izzkTubiWcvEEzkhKRakIbBGeN5cYtUsDc9S48uAvh7
MKy+QjEzHxyyw5oN41O1af8nXGLNWJnhgTKwqahfdzXlnjB0Xp0gk7PEyIgv9vVkef9Dp1WMhUL1
WRtQ6KUFOGEN37CuIX0Dj0n6nAv3BAKVpucDUsl6hyppGfdXJgkLRmDAJox5tL+5014HL2/saHWD
hYonRz9Cf7ea7Y+QNsFS9N447/antt3OYlbA3bis0bs3at66ArOWfU1iunl54hz05Ml84ehhAsYY
jeECjq6g6ENGiVzcM26mqhSr2YGCAtjYi+Uq0GxT03+yzC95kTBPHq1ZQ8guWpLWjJaHYDMSI57l
o+dOtQJYq9ym70Wk132R+XzN9zZ0ELDf6ge/mGPUN4eW/HnqX/WXRML2RoC0BmFdICCkXDhOxugS
61QVFi7e9KbTwgurYVbPqNBwxu0ChSedGJQ8baeXK3hndJmVAStRCBVkQxRwv0zD4GIfgr92L/Ma
5Nvs6dOKfMO+qAh/aSisHigLxsjpOrRj5gfXdk/adqovWb86WWi5FvDKjxzmg/8Eav81wYuVdyuX
c4OuaKpCqvWgl/3dgzyzqCmX4nfXIzaUyItuiYLM9U58rvghZ8x46tIKloju2KSSn5VXwlqwlC4T
6xZLyq2ijmT/nO5taKzui7SxVbe/7mjBRj+XZ8adHI21QfLvZtNhAI7SGw/D08QJMconch5VDwgX
Jbmg31wEJDiPd4b44HM+EiaShitMolS2VQv624slvApdIieQQ+yj01QyGGjjCyrPYmZ2sitxbVCM
vWbnccPmVOI6A/sSu/ktYkrcJF3D+FPHKlNEML4bobrEiuxI/AlP9lYrzr+cR7ymAoXDSsyOdTPr
xei6I8fenfUBdSdnr5PoIMcixLHVyeyelP5/graCWRaNTDOEFUoQSQD52/PgL2DfWRzD0qFFdNdt
IQ7B6gRx/9b6mbn/y8IQZW24BN6UWP9Kvkrmi4ioCpoIRT4f6K50HgjelUGT5QYTLAhif5rBwVu9
XGoVye5XWJnMofxQV70Ank15WugEHRf10YH9B3/P51n8FtorCrl70y03nSzcc/+bQs2OgwZwjSwa
LPCx6dZAL/mj/UzH35f3U9VhFFaURozagw9/CK+j+lrtu8c+hAV/efbDMbk6hibTvt134oLVKVPF
mLMx75KIfgVjSaOBDhZQLyQhn3pzg8RmSCpeZkBrnVDTGxMgWxmmfCj6URz5pvIFdv4zpbxIWoRW
8iffKrHry8ENKuT812/tIga5o8ssLV1eObSrytsLeo3fCHZjUPtwlYh/2i04NHNdXq9N7aZ/Prvx
4LqvAPZpMdQFSf8ixPzYucj9L6OVu9FpjTx3wZ42racSYQ1edOu20cr+d+e16+r7zsDKpgrNHpk/
FMLgkfuEmNdP93zQ2YsfiTpchWYSdWwJXEeEn/sYJJOoO55fVYhl9Bbx+PwinqQheUBJ/6Pfocqx
qxrJofpryr8zMdlo/Gzx442sZtIjOqAERVHnGE6rxPqMfDIINN6rYqdheg3U8gSyLfz1Ym/HUqfN
DPVF8MBHaj+/Z8l5mKiGyQ7UT0oWZ1L6b030vQ3CKY5c7W9ElgbpJVnWOqzdvb9dV3MYZidIViEH
e405p+PxW24M9+mKs1/yKIQKYSvq590NJUbcGxLZSMvAhXpFRlyWm/B6r9ZdD/GFsbTzjjJyTBRF
lHSG6ruWE/LLvXeAG0dGDxMk1fbsHgbPC/RnHCCP+gfPb2SMmD2/rKi9DhTnS8JNBXDYScIfCrUI
OwHYUzzbr9YsDjO2IbcwqIKZTdWBF2z/AZpQZx09XVpkGwXWZJVB7k+kdXxQ8G593W3obiLQlheg
4zki32gR8ZEgxD97Shtod8igM2ac7QgYQAQFUXNod1Wj9Gqchcs2Z54/jJvLCbTOhjUZ2NMdX/84
DoZOpiawHVW8KiIEkskvwbhp+n+0Yc7u41LfMow5Bxzg9XyRkzCbmU99+nJsTGr/NrFBnwjRwfiu
X07f5B9yZ8/DygE40YLENKrIImhNS+K2WCvImy+JVwbdNke7TGcAUQvz9VjU/IbtK1+DgVMGD+lz
ptH3ypldYerJhQQuq+QHoTLJX8Dqlj9GyyCOVCEFUaXkc8BYcybgFlaPajOkSts0ycAriBFsvqw+
g+8ezdkyHj2v8j3w0Zcmi9aIdKJQhkGcaejuRgFvOL6+HlYPZNxbQwgp9oX/m4iBCI0b9keNZAAp
v22aTPQovUuSYvC0E5mUa7TlmxPz9yC8h87x7tbR8XtWyi8+sjssG22NXg986iqql4XVr+lCvvd9
iSzjnnB6F4NhQV3jWu4oQVPR3jCxXCqJfh4jIiLaa0WXKh9ZxdtzqqRbrSpqDMFtmLhuH0GXr0tA
5YLRllAvn3zMPkIUfJYjfIxoQqonF2BkmPy+hR5eBM9XM7Tb0c+5S8NzhcUT0wBTrvT2OxXtDQ4a
w1Ny7HNOA1UjDBGjOcVDgmudQRRR3x1A2EGuG173Su+NTFW//qUhsqrzPX+g7QhNewxE/pURwYn+
vzRbs+KkroJbNPmzgFTTziCQ3fCwFQBWu6gHbwsjwVO96z5UjBybuwLpENyzHBhrXPhuq6yJUY1Y
mHNPezha6jX7JBgxMXN7KnZNecoBjjzXN30mHLu5APH3h8dJWPM5uWhLK58KYEgaf9wZTX5v8kpd
bDUBV/viw6CuaLpGpkieVB0gsF8kJoOHkB31q3dzEfZxy+W2MeVRxkeFIjBSG3bqu0Iy5ZdrmqrN
oyb/XWK10cCwE1oPFy/hfsafO52mYMfLaZ2mwRlq5iWO6DuYh+QMHMgw4NmG8SXWI7SkigwlQdE6
eOn1mUp9ve1VvYDsHef1v2SsEfVG6+CUwBfWGhITm9SDZ0NyKoD5aOlT+CIoI+aGqD52lcz5XLiG
FeSkbmmT5Ho0aIFvWBmoDKu/HUOz8b9EQhAyEEJOp6nViZBRFAv7UQl25rLJfNUSWWS1Z2LCv/YL
rW5/bDr0HW+JRnXhzIu94lBvH4OLN4x8sbY2Uc/P53C/ETWUFe3CZ4+vkYMKuc6qS+10j4yR5mhj
9lHTmxPWxpPnJEtRxFV6cAy7dQGzScAOTmjl1allyHMpUpMdEFe/IqXWaOsrbb8imDnuPR2/StUF
+MffCooin0NtH5xXvV9sAxP37vaJ3ajEk5GQyX3Z9G1g4CGIyWRjLLYCDE2ChLtApmC+59qUN4Ev
m/Y9L0logVMiHKGd9TEv3LHSUtUuxlura6I0ICE9WxNIxpfmNhQX3O1Uc0yn3l1E7tuL20ghN13Y
9uVQpONMzljn24uQwI1q5frpzHfkja9w6EwkOfhOZhUdhahJfjfSQB4jQNwTOhxbRgeXwkYttF5G
UlgmILaLs3/ixu3UbTAQcjmTItufqS5RlCWAgqZoabG1QpUY2psIQpoJpEtZLTC3JMLQ/xddkrPq
6EryRXS7DKqyO4nVtOjtcOoRBlM1rCp1Xi7jTdgkOTCLp3j9f/BK5AdzD6yRq47e8h4jgHhnxO+c
i3XPSrhj3+twuS8Zo0TouBvcZ0X7LUtlJ9iEqQNmH8R1o5P+UsnGMu6V6rRToOmP50al1jfPsHCR
mPhWrI6rBMOTmOWtCLGRvFwGUTgJ9pCuMUmQkD2j9i+O9c+IidPAHyA5jVUYQtAtXkbiEb5Qi77A
1h9pHswT5b2ybwWLcpdCddI93GIJVMiDnn1GlYWlq3N7SWX7OVi0tFKmz2F9ev03GNi2gH9rGHBV
ezegBQjr355Rr24ViW1c0YCSae/Hgvts8v+wah1Ax9PQ4KguNP2Rqn3h6O0k0CmpHhmR1d4o5VVG
5VkAdPlgb8LJEDKQvdmYRpH7/eghLfTwIxakPPZn/HXAZ80sTQX56nQiBF4j90ZIOqTgKtsk6545
SqZEkHfE5LFFZXbBzJSjo8KxxZyzx/E8FJTPtfX/oso/Phcr/n+csK1MhYeT76JpVUq5oox9pBk2
6gX5j5Kn4yPgeN/yJGbBBqCAhChbccNMAcIYqkk6kZlulCNOvOuf0tlI7YrudoJAaP0ybBVozeOR
gJVsNZUpYbqRU5uozFSzGgentYf++3jfdxvuQKUCQFrVUPdkeJxCdsy/cj1QzfXTpphNMRwn//6o
KLGIZ4DIY6foTc5Wt74vP3Mpgxb09IRovOsHmG9dQpalXIVgo+CxfILOqLO/BcAL9FkzZTeAAN9y
8S7IdrPaNaWqHNLy9ipv40JO4maFGpMMhmtodNq5ccpwZTLCVSlqY4qW1VFGU7f1/6RXE9LFYw7p
erTIiRAQsjOKK2WUSb/K3HbxDv6PzCKh76XAgy2ZwYd3sMUe09XIrQJSdefNUo0WekT4K+aGiApp
lom9NDNXavtj76++Lxzj6b4EWJ+6An2VZo3h5zpJyLLrbVH9dySrc8/Rh/dgIAatYQc/NVnsv0cb
7KmA6Figg9MvoQp84naMQVKWFqXslRdOPAwE4Vi4vWxPuDeVPc9OYH3YA++PELYWTw3N7lk4m5wG
h22owdKxBX4vHQ8ykTzrBpSrtmV1kUkdg3Jd7JeM2gmTtgo4cgT15nRkdRqTpOosPS9KaVA8bqdf
RNgW3R1heKi5iXC5z1AV9PvSRDY+LL06U4PcavcM3uM8ZsyZroJTcGgxIBNtcfLeNVvnOvIb6u0L
vAlTmsV6vRKPO7Pl85Ui+yBqMEipLMddsDLyPl3lubfauRenW9lMl/sRijSGQeynZB6ODt9h4dKM
9zVCT8lmmmwDaWo95GaI3S08CIy9Xj/3b/VPoKqN+tdu1JjTChPWgf9L1eGVA8RwFWpiSeY9VGUB
YJm+rxZTlPS4VZOpftpCqCDaauMcxuDwX95guW+/GzLfzxDsXtlvFWujPFoaSy4xc6MpgYQtYYCe
qby+Y4W9AfEkMK5XkcTSZ/AS+Dsc1y468j79J+H3d77Eb78jhh5yBgo9nxKu9BV3aDN3g+ANBcJo
RfpzVM1Wpm96SPoRo9t2VPPhl1vcUDCVc0GEDXv0mEoboGgiVkKOaODIwdEf18vM/NzsBCrS/NO3
+HpilZZ8Fv3Z8XjNmaoaay7kqdisuPAoaiRj1467OXF2ovBgJPyzPbIkU9eZjyza8gvtPdj/1KPq
C6pwC9apXPwNeFbLK2AGX/QBOUwrmmR/lf2gCR0Ji7Ckfnt26d+0BoI1UcArJBlaZ0Ap91fEMWR5
A+fZ6570chZ0+KtYKS1r5/9K+4Mm6c8dgjZAQ4muH0i70ME8ab9RuuqoykxaW/ys5i5uDGMj9sbT
F/d9HnNVpNu2gJWBMWB4ugiWGI/bxg5dZCCNtitXE4FE3ez+5EmqzAA5MGksugXiyx4Vl/nWxCz2
eXgZVZquq65VCFTAHs1CxTNeHLeKGB9W4tNMr/SWBkmxeydfMhtKfj6q5M12sJIu+JACxL4dqptT
f4S7s7DPHFdj1Wx481AW4TRiMN5lAgKsZXrEuyZcLNI+xfZ2kPKX8248ZKerdZyra61m04u9cCIB
FCUfSWE3oispYp4J6SgfImoJFAjLOpX5JHuFETlkAAzusCokVm+RAJfQ4m1lzjNEp9BkLvuG0G30
KlwbMILg1rfUmfFsaXY4hx4y0zbmxhJX1oOZeVbR2acfPh5acDwRJBees6mrAem8WsuvQuGdwUn9
zrgrr9ME3IwW3oUMPS7/aOOTsptoARUIhXqGgZaFjhGxiR+FUpWVntV/KTtvBeHtkNXe30fC7dQm
u7zdSHMhK+WElRgfO7PDYayRUhq57eWYG040yg37MpRVHCcDaEpU9aMpSBCF8kXWcfVNvwXUY/Hf
mExcpwBtYj3mdHPBGJ4EQddnJhI7aESEkkzxD5pDvbS15DeFIyxPbKnTdUagDJ48sWlRMeCBoXG8
N8Jgit96uSxtr/u53460APJ1zBEKX4Ns7i0uim8G9reOEbpy1V/Kbm7Cye3CCcBlOIyMob84uXu/
l0pBmKfdTn/KR+bOFiktQ8wlrgX7XkBV7ukJg1bwl9D5onpzvqSe65mtmTwzPujMt1aOJ6gwv++7
YoXjgw7fSibUc4tNjdyVWddLD9iICUWT1kqjjguTDqg7q8n4H/w9Cf4rijlna4TvsMVO/kE9j4Jp
BUi7drcX5Gv/WtMn+AtycXL4jkuIQEoa17MBcVBc7fzOPNHwSzeRHPKCZlV4IIp2fJ82XYZ8dNMZ
/QNhyTrOJw9rTXAlC9P2k4Jrgk6vJ6JTKJfwM6yZX7K/yDWfu3/MxmpW0K0PzDPuXEPDm6VNelaw
KoaE+UIwMQZIbTSgEmXA5L4+CzjTJzP8Xh5JdX52RQ+8pk2gP7XRRxFY+zUZiy5JFkj4YO27Jnsf
yMFa9LpwwtwFpkA2oNOCs31kU7J4L833zYbsLCspOI3vov3CgxNSYe1oevZeJx6VY5YJwGo1P4hn
elKkcSV7fXIEnzpFrf2MPxcWXzlMUsszeOwHA+ytB8I1N1XHZSRu6rn9vvQDtn2ok/7YwznGpWtQ
X0xYc2Q9xNhN88foC2VVTauytrFcNeptlvx5nXklQ+kfPpqnif9ujcEnj54VxHPtHJIOI//+vSDu
E+57oWzIRuvdBGRfH7FIxp5Wq7IJroQRd6Cxy2ual6fw+ZUxbyiEIhkXte8vsFsWoclKZG+uKrhr
DG/j+2iGpyemNtL+0sWkPdC4o89qMOR7tVo4r9ECQsGyrwg0AlsAKOivvQ5/K+WHH7E7IqTPEEXs
LlhVBAPQ3aLiKPqx68nlSrB3+GlJ8/XUlr8TO7hTGFnSYO072xh/kNbFAIFnZH7KtR7U9rlnt9Oh
nEzd090opDTSWg6Aqyee2zOLHSnoifyzOMikWfCspNNO+pewEI2/qmb/O9xtpBso0k2R2qM8ue3n
fPO3aD/e4gF9YASCnnOhygALUCLm+1THVQjGdL8HRoGysI90cFOXuGU/dXhPob3yRl6ilxJRXzUO
SiY80PjBDOYvr6whu0nv2DUa8boFfeeMHdQH7veQ/+ZxwluFeWOLzNCKJouSwlHcs5fPavj62xtP
B2pQbr5PJ1myYnxBYOlIo1QJybis4npH5BC8zMcen+k4rjIAjzGQrOwFcQJKelHsEXRVS5hk0yEG
eh1rQf3qfu8FJkDD7cJehNAmCyzGEVzesv0G/CJ4PbkYZ4xWoOLDv/9Dlngx9MAd4a8Ebb85CH0p
1I0ENvfjvIf8cQ2kHAsApNJ5yHuP+RdNAr8MpkBOXNF6DU1YnBubpuhnCp2s5kO9CrlAS5tZBuPA
jaqBioyhNwGpv9hRlCXenKqWmBMAgVtBcUDG5W4WqS3KoUaSvw8sau3kMDAW55GM0aPYRTzHDmDJ
M1viQ5VldL/c7npRIOxSibh0rBcB7TJ2SurC5UGMX/czNT4hDXkZOO8IA+JGucGdXiiXz699L9sc
wes4TSU4a+Bo7wI+uAA2Y0P5GK9MVKUt3Y4tqXt+yneLXTwKYVYQx+ba+EVykiBUH8ODhUEoiDjs
vFN6p09D22KqfbnSmo24i5qK0Fsv07p7633jaTA1XToE/sykLmn8pssCDmetH8ECrWy6qcZCekqv
Xz/GEA1ZgCmMxPw9hqCvqhE+L7P5a3CkjkQOrPdJKijTMosJdpMCqCVy/nA36c4bHQuQiQpwbeef
CxN7c1lNJinyY5wwqnCC6ahg2ZDU7h9IrYD9fYFuLcrPrtUio6/mt5k/Hdgr2cRHiTQId36YjzT/
/fvuDXGKGDWK4KsORU0irw2IwhciAP0guQd5T6ZFusKxmfge8yy5n46xsGM04vETrSvxFQeKUP8L
lBz4UM+dO8Lrei1paBReElLVe56PD4v5Vkv+wyBx8pwq2DurnuzGWoe+enZnMzBM7TOxayXwjGSh
dh24AbUiBhHFbP55oSVkWnwHxjKSgcbyuF23C2Y23jfprATclabgCoB2EoilKhDmfo2YWbc2RL1l
MeQGExXgG1TyDIxkcXLv7r6DDL4qiDw0J2+5K8XtSWw71hKKgym2a98ytUDNGorIfiU/+4Zg86is
oUSwQ83M5KDRkYpB2VpJuIoXC4KT20k7jR/TFpew68oBAsl7kz57ZrPiQO0oQAbnlToN/HaDMjin
6WU/1K/tcpfH8eP0j6VybqC/MgTbVMTBxlTp2MGfzM0h63qT9r8wXq+k0mfDpPZ2vNpg/HmKPn4G
0oOpyNYZTC9e4zhjTJen6PJjrdiLvHT5QGijMKs3VVr+AxFydI4jvbAB80yp8qMGsFZ/RcW1rbCy
c+6bgX8J6esS3zAu8pMK51TIl/2J6j/r7QwsJCJZaGhm9N4pRrzqi+kjlZRv/sGfRdH4SBIa9k7e
c7l6G1G9eZzG9/ewo37P6y627JLYIPzfKhYN//riXgVCYwMLTN3ejsGr5mQoLnuLlwgEMhpkHos2
QEXGP+/Dq90D5lgJVXmib/g+1UJU9GKmSEI74hQcQc0kgN7+ZfXvw7OEu6wY3JnY6Kuy5OLFKoqs
q5QB0dz2vPGDgnEpM5Ojb9hPxrpnz+B6O+PL0u8cpsFOvHm4Yj+8DhyKhTAWNxPN5humHckVseJk
UNBCDO8EU+SrslFVsWIgVFWdlKgCcu3ANB0kRB/T8xKpazykwHMHrenFmNiArsyLL6mIS+lfpNST
kST1dB9U/NUHLMg+nswiLZ1Q3eiieIDXWK1k2urNkDBd2/N9zbgQh8OJ0EdEp7QTB9RNtZIqm+m7
krKZqWAGjDgiR95K8B1+3x3whywoVASSUyuLOYxE62pyW2w9knIzf4BlskuGAui5PXQApd8WRWYh
aH8FoPbZYzQSxJSp/EjX+ypN8q/vtUh2pup3DZt3wFUCI3AzjZcKQ0pYl35/0PbONFrgnvXobMX7
C56iMguhLJOTEs2K6kjmkPRNt+15YraRD1Porr1yIZgDxsxwDU/Qsrm84aa6cFcl83DHooWKJ1QM
XMOn4EIYEUT5guEr773UzS/UYCVpr531TZ+n+cSv4XUu0xTneCnOij8WwHffMR4JhrVkj3Z8eLA+
x0554vpiiBLwh0LDkWD7eIj2VS1Kg4rIjfMJYuDKCTRzEV2Z6IvaqqAdwjoUtQn8Sto9WDt4mbQ+
2oMMdz8iEmb7+J8yx7zdhlRm5ZI67eWEM/7JlVlfVENk9KF0HDb4KaPVD5VhltpRz4ucY/h/TTny
TkmrVfaOFaBZSj24cEufxKl2JtD4T1vOsl0Ld8hS2KA5vIscSM0tIlmavnL+58BMAS8isJAqLXDf
zPSE4SSvuGkvPX3CY8PFtTIvvL7WQschyy7L1XySe0fJ719FpNdhcfP54beZsYcCNOkKEhrSuegN
5ODVCWldhkX1P+dxoLSJVqiosbrNlrQTKu0HU1sIqTMou6MHY6If0L41UyEhRrE6Kn/s7/5Y+qTF
JasA9o/OJ6xZrdX3A9j4/BY9zPH2erIgwaGrfZtv6+dYAU+HFOiAXQTKCaz3Rg+c0xZBcSMyMPvi
FeC32BzVq4bTenRUlVnA0dscRI6MdPmsSKR9DCsUcdkVOnTb96G3c7MZZVuWZ2SGRH3Ju8yWuLEd
rCzjU429KnTxitzDwt6tHY65qFFL5aqWNa+U3FOQd1TIgCHLLrg9AS3j40r2D8RJU1HQPg7UYSGp
LxTNLKXFq0gM8FSqMtr8BMXbvv10rahQVz7i3Y2mAaqFfc1nK1+a7AIBPrcnQcoG3N/N0i1ln4AU
a7ePLsn8IkmEW5mekENEJ71/0MvWFsDgQQHeGODbVSYXBJ2LGFQHHcU9Yz2Qjv898AhLs7P0K301
Vh3OrtGgMt1Yb1FXXaHG8ByJ6W09+9EvxPQrK8DnheMUtHLo+ebS/5PZrVjUb5tyYkSKC8labr2E
X6GTo6PHyXbaskMq70bblEz1A6g13emKJ+tD1O+fovnLUcrYBtpF8+EFRS1zRrQoHAopdu3NCZsM
Ti+Ug6aAPjEwD8eklnstLK8aYTTKqoQyjXcm8YB5dXzAZNzHTc89mD8jvsww4EHVQ546UxdH3jeu
fmdqXNRsWDeU46pyaRSQ5I/bEhGCg4pjnU6ma+udlC4E79WzMejZh1iV4VIwkL8Db0Dwa7hwFJvJ
GjR36m6cSU9ZTT1j07jgiYH/CnXgqapusfjTWMJcoTdlbGqsZUKBH3gR68x5q4lMt2+xG35q2zdD
yYHPWR7Il/oIhU4YRUUN+fEeNPoZkMe1CmlPuOS+dImWG4answNAQlSDrSyaZug150m7LE4PYmwo
WCd7D3tNZ24jCderXiBre/bnRGjxdTukc0/k0ev0i1akxjmgkHQFk1TDRljT1i9mwNf2h1SvA8rD
G4XzgBJSH4PPSJt/Kj5Vl5Kajpba94mS9eGZeTqavY2hcLWNciQZMIejhavndnmom4SBGgnBaHPb
sUvNV/dVeHgSWtHq6PXWjUoWCbZ+ZVfbR/DLaivfqFyF5UIQeSnjAvOXeOfHJ69O4+LPBN736FyW
5bZCBECbwgKLk8A54D+48Xmu6nNzAKjFU+IYs0KvIG2G7PjDEJo2Ig4H51KsF/c+OSBMCaE4VwpB
//Lk7WwfwzXuqBMeayiiWY9G92tIBT/3nGjqQLIzjSXyuPlo40NOpPRrKrYswGVk669L1I7zps6R
u5qfvpH2PMW+t8SJA1urwKsFY+g9NFsj3FISq1dhCkZaYp5MwXbH2noO72EcTmLUO3RbGcPreUlU
MqzDE8Vfq2WpXN0rvd9wCfjHrTlDzCexy8eoq/v0CIWPIa5I9Kvy5u9W/omZmzPnOi4vYHWw3194
+FIVSyMuoERQvxDhFZqRNi7kH0J3z4Mge6iMr/jc4QhLQdqX0RWKEyuML5Q5TgM7Yr4+PZ7in7bY
QLijK/bstBxmbP14dp7O6p8dejnIbU8cbv5L8bWwtqSO3cTpb+3TQC8Yotgh/T3qq5pdjHNp0Ghu
EdYEaWpuRpJkbza9cSv9ONRwJkrAh30LahzCMtHfXkYGmF4E5fXPXlvDaRzL9MZtqmmX/I1bCE8z
TOlqdp8rIvStu+Q2qra3StEnCZ0uS/1LKVSCLR8gEFlWC26vQ+D8CXMklBboitDckGyw/yu5xgX/
CbTTfA6DEA/rJEtNvsJuugEoIuueVcaqLlhUeneAyA12jmstpk/d2+C2JEvOnHOPdkBxAUTxGb0X
9BXzWy/XyNWLgu7UIqZ/qpdu9Jsk28CNg8YlO3a7PKqG/WjgTK0tZAURoQX+bXPcRu6r5aY3bm6U
/obXLT6Lub6DZwmU67eg1Q8xl7WBGz9GSEcb8HuNEvrsr4oShPrygoh8wfBrhOBLSp9o0ESdFs2F
W6tM2PGJrj+2TCbcgGUA6egaQecNhj1feX99aYmIRgZ2Bm7x/jmsnOBjEopzIuHtwMHSrO4ep8Fl
UkrIfwti6bxNqIh4Mn4oSjuULZWdUk5pQtalMrtMp2BrWeo4j76VUTgTxIKsboh9/q4PSKXr4uxA
EHykw1Cxq5MGYRYsaQ5OaD9u4tUmjunysH8x0CQUb5XmBD5TZegy2YzyVfo7NYkyzva0zI+PBk8L
9Z2R9H2jVx/HHf9wxCFgmUsEBCK0z+DohTqMjpOy/V6NBdCUjXwvu1J4U/i/jVYtDDJ+eUoPANuw
SW2vLXwxF6XQuOp+fdRsfsNoYiIIsDaN9JOkQT3fy1HUjP/KjmfVbn06wpwJwTiRYa+fzjDBtuBG
fld/k150IyhmvBh6VNjgoA45OWe2mhYtG2G+5txC/ocYq203Td0fLuj/LC5gHKypCAaWcJJNd4hg
FOf3xxR/UT/nltxHhAWTxKiN79hyEplCNCQTKetYoog0yt5gccywXHrt8Ruu1q623eduABWiAXmL
fbFyZ6rtMAPAGY3Z0BimyjBeoNsVxB7UM5nz8bxOv+1hVi8NGW9Bvy4+VBMD+gjBsHqI9XEA8KdF
Ap70pLDjf0yitVYUiQ+h6g0bEecV9MO2A0rxSeGzauXrqoj/EhxNOcUqz7+13BxNkATKw+BaZtyn
MSkmcQzCwDZpHe4pyiHAcvcwfkCoDLRMPtUzFf+yaVzNtmdN0eev0kCh6RKYiHaudq+ONRuNw6qM
fFGcBy5stg2eKrbw5xXYWxayg8asOV0HCQ40/RCRWS3KNhs/MKJ5njYhbraqaZjbyFw3fVB/+3c4
iu6aZ/dKmlt7UGA3Vqf6Vp+Fg33Yn+Tu+aVBQaeeRdmMNK2pdSU2j7Viq5c/XyleMF843GTkiYV5
luJwpmrs3Bw2WHyEwQ0QIURRlax7rcZ9ZN+FPPrK2oAG2GuzYLcpEaVufRvyQZiKm88uSSkw73N9
YTvbt7kGml2npjqkvmcYsezKEzpey6FHYHGYzzdLbdeYUZH8oSIcLoMgvFPwHJtq5sQ6SymqExv5
01SLHGRKndsJKJtlXXUsOWOpcDw5j1ADqZ2OFFkjOyZ9QPqGNBKl6HvLHjmcAX8dYgtZlBs4U2eP
FfRfCe/ULVi8h++O22WwyMGzSgWQsBuW05m7yojIZj5BjNN48eEkjnZZ0IeyM+U/sd3+ltgvtAXI
l74MTWaWP5aGLa7rCObTFF70qdjJWRc4O7xwSa7jelYRrVs+y5QIfpHtk/gTdgPw7RQBHn9UJyEG
AuhjFMFYVqq5tVdg+6dZ+UtLKpHLVY4lnKMgBckgl6/pQSdGTM0TZUspB/5rA47m/WmmGlJj7P0p
0yi8GjMd9q5867nQM3ZIPw203LJpw/4x3rCG534io5oAzqnlxBPVlVm0qC2woOFzMgMj76Znfhr5
fiTj3RCdtgJsj19b52WFKPoqaJJhgIe6hWe0Bb/Svzz4NFjU10vu1SY/ruHL3cHKGD+rjSjkti9t
JKRnoP1wB/qrCIggeeqfdX9wGqEBZ9L4ldnS1E/rYf95MSndAIgyXs+pOXgOqucZQOo5jYqjhYjj
edRAR8R/C/lGeJefb4JdWFZWAxLTB2XQN+52y3EMFwJ60iptawmNSv9I4WkV3drTN/uSRODzM6TD
bOohHhEGCQboQGy8q6GWvaYSWtEULxe+ktL6/H/i1PLR8BwMeGNRJr2prH+QGSj6a3YQBBt9ilzi
erG9sJLgEILTBRgtNUeMNxa+NikjaGb7OGCG1gc73gukpBe2BLkp38vAXEJ/wsgnqUF3FEaSqtEI
SqZLBDmljTlVQu4xadol+VIrFBF4UAnLHkEXjA6Ny6km55Yhx/O+Oiusbbg9Urq/xvtpV4BzF6s0
ziufiTAJKpCKljU75QieJvv5Lp/aNN0RWzWg/lwAeZeLSMVz6AYxUnsr728cFz8Tw5ulxrzPbc/J
5isPMCDxYc0SvJCwdp+qAkrHJmRhqSFJHILqc9MVycWiE1r2MJJ6e1xe/HcEynhh1I3Ur2hVvWdq
j9lM9oIWwU/Vt3zuwvS395eiXs8T4B+i07gdRvCoVaSjrCVco0431Wd0ACqBUwSURtWlcY/pRhOM
MIdVboN3oGUCwhqsQ6NiS6INCaP+gzZMQI2gzU/r+aHKFSbwtlHZ1zUu71/e/eLjsBbctnkLZxOz
BWdW+BNbidovmNGmFwVwcw0nD4/tYul8R3foWgcBL4kEcq1zOeIyFUsXHxLSzPs7Bgi8EWBNKeeO
k7xVGzi86ZAmz958yrldH0dKxkld8q8ogiffnpvMXAzu/5XyWhBKv+XNPi0IiUPo4eVlwDtBfhi/
Yr94QnGxghCFVRJt1l/v93vv3Yvsm1QfGZ276T08A3EMCEXfzY38yx8bDS+lzCYRRKDP6Ohz0Bss
1TRZg2cvEina9kYTsoZElRBKXDUxPBF4onMde4dSj4wlLaVEpWOxG3mVGGhGcv8YMjn+RUx73Y0r
djv+ipWfahD44luSS5XCRlSQzZxTke8aXpMaOpSfFhZK3WJz3rJI9zN5c3VIS0pOJOvYtV/OHyvy
k2dtH64WAJrlZ5j8RBZoAnsv9d3aruUpS7sZRmK/74qkhgZ11qWGjoiKb4+a84+ru3IkQjPrmNhd
xrHoUE0yIDp9QRrspfp8+91ax2J0LIduDZbcxyjyQkGd/Hip8d1Vywg+/ZCZmv4zEpglDBEJqzWc
/vA42l1J0MGPEroIkGO+HleWOhQknGh00n++BGbPDvEGga9xNn8PO0TAyv3Zg574cJbBbkxRYHgM
fFJly6+Gxi/qfst8624joobmoAMWn6vA+rFeq/6SS5p27hlXn8tPu37XGio5MavYIzKovWR3VURF
LSOw2Y122jhQePTls7S9QG+ZLZuLVd18gMABTlp2vT2kfKseId1U0QpHYS0C2K5l6wt71P1Irq5b
oS980+wVaaLB+NYx99zIUNhQ8htvhQrYNa5/DTdo3Rrv3YnPN68xOaLL/XqBaFY3az9fhZ01ZJX7
xgFYR3wgiCUqA5Rvm4s7YCPBwiz6BlqPhmglAfRMqbFboWwaPusgU4SJpikLaJnXNJtgPLCqpxVc
r0rE7SZuuig1Gy15mD1jFjmT4TT79XO9nNnfqmVW4oePxXr48SyxCh4TZS9rJXv6Ap4BBPTtfDR7
uvyuDMjaM82VCqNerAr5ivksWaivHdNZq44ey2aWS7iO00vJfSBeKNSeLODta3eut9ZzoweWNo7R
FLbSCzlsxse/qklgTuSQ4BXIEjNvl+xsdwR6SSMfD9GFouewysDpg3JkXkSM7/s9tkoQcY8yFKvz
xX2r01Nk0dDZYcEmXnydNqVwO8KFf22C/Q7taIIMjr+CwSkABgDl2Q7qZelNLSPRTVcWlaX+/PF3
vQOFwDG2PD9ju+lyCspk2i5wAiNKtbq1butNgVSrCHI3w47PGfq5r9d/+DrC41JdXkmrInetwDqx
uyV9uwyZiolaF2oFmziZRj2u/OZidBzvUf+e+wrPfZmiNL1xk51S0hLxtQu+g9kTU8hwqzlQ/D3o
GiB2H71qH4/IefQ0W6Ka3a0FpMAOEmBPW9sMwuWpohidNDXSCUCd/iHTTC6FAMv8CtLRf5clXhcD
zmeG9LZQqD9XKKJBDdysbNIG02yAdv/Wd/djkoa24OVLGaTr4WIWeieDNrKevdyZ/70W2O2XsxYc
LbbQL4buvSsukMKu0YLMhVhMLhy4LkCTMON9sKz66Tfiz6PS1kKTf3lMHZTDVCxra8rcHhhTe3dj
vP8BjJuh6aHCEsNvV72B04/6Skzj065hKgF+vHPrTRkf+V9VEz1LS95m1/EKdq6MDgIt2ZbW9cij
hpIvlVxIGAD0pjdrtjDr7EhHiw7fTmfzd6aBB8NcPbO52pqJ8QIZFSc40/cGJKEep6NcmWqwUR3C
tyAiLlwuL/X4cM5+o+O0aJaZDqae3/25+WLboxe0y1bUiiRzR0rusc8I0He526Ox0S05B7deqVS6
ATLr89bSL5jD3HY00fmMBrz5QoZPbrJ4PGuDEYkGrEtCkx6hoJHcjggDKMiMJ2tuavgqvYTMyjqs
WXR5ue3ejF6giLDSwELP1xvq/6lKwjubCYfzF/g7rWLFdN0avXL/T8WfviJv0AWmeC280dRfS7H4
yLzGMz/d0VDZVx+Ecbqi0YZcO3wp9t9CMyZ/Z0ulZo1cGHQ3FepLpkgQI7nugWElHBvhiaQIgSM2
PrUVkMc2zC67YX3uTHxDiY2Zpx9nbJiDudv9t3jzma/WYKHVuH1RWT83i/qFs4VvAZxBxHe+YIDn
nTWXIGoEgj1ZhWF9+Fawm+wBk54gFVOZp0rv8b7H3/BdDJvMp5AMPbRNg+704Iw+bRTwCDGZ9F5j
CohEQmoAaRWwZB2wFWZOhNJMTsDKtCN+VNpBVsuvx5+DF2DbBRAAuyRf3cuO2k/xHJpwB6zjwtZt
KqKXUGhMbSPOkzBC36NxemQ6jXxix/ksW3woBJt6tnc88aTaE4/dB6akXlHGekPREgHSV1Fp3jr0
cNFint1v4IGZ6Wk4jztGtHuX7qcx07p1s/1A2KaI1XqjsC33ZlmousFXKB6bPAyuqjLv39RShwPb
U/0/MIPPREKmx4K1yOExiHn9Xp4d0Wif4Ej1OO5H3GRqqK+3d5trAX8AfpKdm7eR7pYCX3f1Ns8n
H+YhNLXe5vvmdzZareSa4SYFWuJmLG6GmLeYOMScKUIH4/encKgXgzWHCQOAE9CDhkbpUkQ32cls
Yok1B7gQjtoPq9kvBPHFdDVlNtzL2mWsoGk8IvubvnFJZn6EhWzO9sdiaAncsAoa4P5qN0Rc7O8s
jnwKyAOJOjQCHQ8xC+dJw9LvZBaeCG0iW5bQTYPHijTJZQm1/K1ngDow9ab471955Ey7xE5u0AYa
HPfI8CzJ64eSt1S282x3hftAvXNMbOnPvWrMEXaq3ie0j2G7GdgTfRtC/2w9nnDikHbsAcJRRT8e
RFb+anEdT4mMLqJR6635TtCAn7GAoLh3r815PDU1tFGRYJ85oUmcNWqb+Vn0NU4d8ZK4b+eCkja+
VgEdXgYtF3ldDnXoxafyrxk9E/Q4X064fvxdByXZUiHgsyMgAn1XkzJN/gqt6QD/y309hNRbKgz1
0uzRLZgTUDmfiPZUQLUzauEHGRkgmC7Gk6c54mMzO7MKSP07bvbbKdjyMpDohftmcwE6t6S0ra0J
aEbrnfbEonBHv9KCK7iOO762AGMD3v2eRvSZLs2e1MxVwtbyRF5Hx/zL7lwiINOsaREoEAbAqyfZ
FE9CvlBkZiYJ3qCBTt2LqafTp8mG82O0+DACIApyw+TSh5wZ2MEZHoBl/jhAtZq/jWVezp3MZLr3
DAKvxfazgm2WW1nrq6ndowwSIGsIAtOGkfffVyJXRPe0OXdRMcMumG8YNKV5oVfxkHtdQjN/du0y
KAR6ezCf+w/2S/Y7GDAxP29Gc4kTiDDYhqFLW9fvo9Ug41Gtq+s9WvQI+7nhDiXB9Y1zCGVBUgiL
H1QPpmI+PqfMSMCYy9Gaua0Dvyb0nQ2Uk4VNvqG2dLwmY/aFPH9k2qi3zyOCKUszvDydMo5vOyYp
+OjjJ7Vnf3jlVrdGZzV1zI9dGFvbY7JSjWMwkcsIlG1C8eYuK5kWKZMkS0BYuM4uoYn2SwVt+Z81
osaYwxo6NAdFzwfUHD9tofpL+DApgK/pw5h/gADm2txiuDgqfhvY4iJmIxFKf4qmdNjuOjynvLg+
hug6A0nig8HLUvap5zyKhHwo2pMII+KN+KZEOtE9kS59/EBwEsEdwpjiG2tjweEMGyg1vat+rIQk
Pe6dzw0sHXpeheGESI1PFd3YJAk4PrlhHng9QN1nPAc33Ojvj3zBHEN6n058i2mZDpWCa9qLFdZk
/8KaBjmqQOBkA5EtSqhKn00y3AEG0eeDmM5gprPJrqFeFnAoJvGjbER0Ke8Z66TuOBi4JANzaD60
Vc2bjnEMdYxgfU3tFlSUSDnb7t4JlEpwVYXvKWUVx4lCLh6Dvjl8lq/A5D/wilKos8ra0m78s+f+
pSHQv1KRnu7Z2vSdhe4YnqxZRPqQQGDmDOmd/R12xY3LnrnODZxf+l14Xv9qharhRxifLJMgUgdJ
yv49ryNBvyZFYWSIZvLiXT76FyCsezulVgA/wSWuuLX3sSSY6kJ7viGSE7JLxTS7g0nHw6LcccUJ
r8yddMc3zZqfkZElrlFYFgLdyOqL1x0Uv00lmkZEZciH8/lwBRys7A4vpQJ71/iU2I3rgjyMKNCV
kh6hQ0M8yMFXkhvf16+93PtqpKiEB7x/F4v7hF3Wvko0jLP2xZWiTB1VqeA0zUaQlci/xvjpPLsm
RLwEHSucgNFP2/+CKb8CNbyPR1Oby09IIzAdV4x0VbzWn9eFswRL8VXSalEoFTxOIqW8ZJtsiEzm
zLLsWWAsNuvQ4Fv+I0ZAA0Q2VrxRmEnrWl2w7IMRVOJhBw+3Dkq9mPsTqSfZi29/2kKvI4LKCRRW
q7QkyIND3aBaZDtya3pwC33JwTxPiwDI0Fan6tCyaDhRB9v6+YReolBjalgnyz+8ftwrlheW9T5m
U2I/pv8fOFDamxGD62vQDQftybAQ3jtoOhzpYz+UrZ1F3nZ8y/PpstRYJRlSMAr9CjaYx32b8/Xy
ijMl1Q5H/8NalDxvIoHkt1ef7l0mGSTqJcKg2aa6Fc3q+UW1X+kOQA3fVo7IFlhpoerky2gnUxEV
0Ks5Gvbuyms7vIQIRptvfEgtSgDnhaP3aK7FpGRTIrKQhyQ3hoKa+AobzlPVJ3lTUqeRFA1DYBJ0
6FlxfU3JUZV0e90L6HVc9h3ey/ySC4L2A6xBO8WZBr4os3xJxQ6aixl0K+W7Dei8bFe0d59jmC0i
bf3Xg6c7uF+RctZU+Lk9BRaeUREXLPdgCZUxIrAx/mnsKptkRayZayrsRscb0fIn/9ZdgOPntp3T
t5huMXLAo8lM0n1UJkb8KB5Jjtzzu0Hm68gUY9OIpDBnGj39ObEAD+MoJ/73gpIT4UjkLt8KUrDF
KcmSC1d67dUSYC+9fuqedKqp85yLULQ5a78hCv2WNQXit5znKP+yeSD7b3EGdo3RdLRrpfKUBjsC
SF8vJTmKtMriPcarxc4VgxG9Q68RTJkJOJwu/r4E2YR+B6kSaGlplNht8IqhPU2jHF8mY+dbUJiK
WGonnXMcCM3GhbTq1L8vGW2+/qHharUJoCQYVcoqsF9d4mCTMaIXKGgGRz9PKIvXjiA6Ofg3cXGH
wEMI2OGpp7jdQ1ZIfyCrnnT1TOPwFK/VJ5bYrnzJcJOKSYcgU6idGPdz0y9xfKwABo4Yz/ovkWLS
f0pl6RAmJlYxVifPrSuW5MQNbkJPIfsMR2SXUZsTwcnq3wDdIBIfaNpa1QvUw5QgvITDrcVGEETj
RlFStUJ7zEoIqAvs3+N4ltDpJm+NVQDczchYKohhwo1TEBeQ0ovIb0IvE+8S2+/JnvdA2s4LMwZB
5ktl2t/M+HjPJPZ0RSWhuhj03jDkbjTdluXXn88MNzZkzKo20Zbxq/TVMvjbdrG8nbCfb7ngpkeq
FExjI4l2QWMA3KXAIyfew1kTNCnlFcP1iR2fu8RPkSSCGc1rrkGhVnFcrjboHPTLfkJVwfCHmeCW
2Lsrc77tCYFpdJqtQGWkkCP0qh6sepd8nOYfz7Zkuo1Fyqqsefsygeoabd3pTAXF2tkg2mqJBexD
Kn1UOwngcr3hPoJWm2Z5/mBbMaBaMiIWDYL9WFDgHXuVi8TSokyZ2/0zWyUbcWp0Z7LEYBDJjOAv
jEIZY8QERg931VSYuucs8M0x5YBFASk2nO7xEStvKzdlvh5m2Lb2Sic36M6jF2rEqkCnwQ7iW2qe
18IOixrOGnSUxqvMpXRNWhpQpgd4fuO1hoiaAxS8pM/M3jq3xr9z11mKrKr/uXeOOPPF1zC/grf7
RABcZsrdH41rP0zHfaLJweSUhI70dztZzh7q4eksmGeMImqQcs6WdeIsYuHu+lSNjSJsK146w/jO
3MWSdpQyg9PMLFpW7mok5Db10PNOm0aVhdew5ZfBnf8eVygztjvMz86tC9IRxUbnhD4+qv/8CgxJ
0XY9RY9+cm6tHzVXFym0psnahJBNXVpyvThH2BZpadAoppH6cf8mUffHr4Gl6FDCVbCBeETWk5Q4
pFsby0QgdBIkMK5YBuF8g/897ukwTvRbBev0RS/zNE9uKSNi6ETxtYMSpLKpcJkaXKEefjCjZR3u
U/4u78x8+1s2TDEGU8CzUQwN9il2hzA/fp15/eqRERQNWEibSoceF4GDBqgxxyHlh1Zgc2wE4qdu
9NY/1yJZl49aY2Y6N8tPVzZRfH5r8rZ8RQOdbxlQ70uJ5bWfZTuMA+RAifF9W8eWknr53/jQjO6E
OGyQw+T6VTed+k0F9MdUXTyfy4OGpxYxF0V7oyM2Z8jBuo0+vJGblWay6QleFgGC0+IGYhvWjJ39
f5gfME58vksXRDBoOh/vw/AvZXULoU79PMscpfVU9KXfa1Mg1BA7hVgMoLd4lg+qSCk1Gd8xaI/Z
4ojUkPtHovWWfUFgBqWk5rR0ypLro4mQOgVRpBLiWI9oO2XYx0/5WHRHfuV2L8ibDLumYSfzXy44
N6i9xN2lQEanVgN0tg1vQo25xGzjZ500MLJDp71EdMFUfafafCpwvI6WwEg4dqwwGcwHwkrokYH4
KSLymYm3ZSMhF8Zf6R8qxA/xcuUUwqvvUU8r3iShpj1ogYdyQ6CeedgDsl7D3PvXINAV61QJ7iI+
5euJbZZH6ZJksbYXDyBQs6KeEaMGOUX+2UhuhsQAAN1q5DWIWsFNQsknc9ZcoThpSALUHRVLwwEO
AKlPtAOEVqUIwZQ5tzCS40dbWdOuvs63Vp8UngMXeI+6IOPXgbpSNznDOZ734XB5pzZ+jWmhozHV
P3LdsIMa8k5k2nLwDKsXyU0M7o6+CVcqa/2XiZ7u5LBvWNZ2/3HtuadcsDrijj7Uh86T5EK9ca0P
0Re6R+VMAl6KRHLmGkG8EpMHnnLKG8s4bEc/4OPlU5VcPEhN2Fm/x1TLKAtXVKzBGKlYBHdTh1op
XkoVia9l0CULfihoYByKXBz9aFNIAjdwiYei8T5AN8i0a2Sz9vrPm5Uxj3F7uIYM/g/tMP/AmLHP
J66FMGrKUSzOglCcLVVPVbAQThPBssEovs+ulKhv0qjChhgAeePZ6tdRm1kIvOCr9WgKy35aihNj
6lroEgCLgnN5pGBdNtu9Cn7b5pfGJIEIImPOb/cUiqPVhr65LBNZk35wd0qCcJSYL/EEe8NjRP8r
koCy3vr7O6BxwmKUWOh/wKZ6pgeHdaDRCvN/WTOl1ed1sym8abM5LNZel5r1KXTGYWTu5cIZj79W
/9wtrUY0qHGd7poGxiPjLB2Vdj6cLPjRZxg7dnI43yn5Uq++zFZZRXKwNIhAiNHVzd5PF5Dj9YoB
bxLd1aGh65yezEMeH3X0oaRx/p49pYQezG2o3s76SqvGyxgkbVNt8Hv7ZX16If3CYVr7scXwgRYB
i+pN8fqBdYKqaai+lFFFT6r5937BCqC/5MTokoFtMqvW0A1zqmY5WmeRboQzoSNn+j6tsvSjvOjQ
UarLUknbniy01+X74B6zWq6vYpoCzrgmii90bX/xROJYbuHxd8kzCn5Nkbs1S4+4rmwasMwyR60C
hhXAaCdHI0XlQtpcGL+u1ThFzyunqNcVw7fr5GPu7e83yewazEpE1pdUpDMbZARqEGYnsjkM25qm
yX9IMnkKewtvnS/sQQGYp9aTUVbvX2Q15CW9IGVygE62tlU2TBBf5HrpfdBBrVJ+ghx7U1FRdjCN
R/PkGfUg/Mcn+PKY09S0uoujdkwjvDQLEDRwgNRcq7X0lrU1KCI6YSvUjre+FvHIGCclwXmhZe6T
a90wD44/2smtUfyChu07eJjx9tTptih98XNaFWWoRrd3pZcEMxuV87DAF//3mY13M+zFg1jQlPYI
sBVRT06jMwUUx9AnKLDxH2Pm9BO9BzBTe2oiVby1KK6v7V0PQqFDqkfc0xF4bv1VtBIyP/2tGFI/
JzH74yy4nBoQOxFJWLo2DCwh+RqAgDvOAJe7bF1wJTw1i1bSPvtlg5Bdl+ll8YPtgLehnRtb3tuf
NOXBVv/tx5aDXsxTS1DNlUHiCNKsFrwsgnozRKrpDPi03gwYqVHOR/C5fs1tUG805zpJIzTho/FX
LMv9o2LvQMpO/TbZ5BIfOr4HjQFRk2/uPmdt3b8v904so40mrKOPEIuZ6ATp0O19b57o69YIbmF2
YuJ8oBnPESuuoU6NBp4UJNw821zPuWdFteRDf5aZwW5T19PM+4lGfilbDPAhawy5GYltwPX+DMNf
s29auZGzM5kiBCKH4xjIitpRrroGWEZbOKtEAEGNJE6rMtHv1+v5BTpgknjE0T+7YzYrZFmH7bwE
REEy3tAU2OayszapPNKlio3JOqaOmh5yUH4nOCSvYszZ7UEkaNNXEpYce62CBKhFMuQi3dnfC8Nr
bVGcevIT0xNVoOQ4TWMYLAOXoA03wJaynPQPnxokJbwUZkNx8FJBsNh4CI822M5eXtau8IvbRABT
viFJ6bT5ZvL9D90sHuzaELHUzK6kONbyLIx7AgPP7jCRGfl8WY9HXi1kKtMVjTadeJB/rDSAB0mh
ijjU7Nmzjd4bU96LAjJ+g50qITkm2c3m/fvjYMphzEPuNGDNTMOj6NA0UVh5uR7CrQfxz2QKlLI9
2DfVjrTLPYmypTqC46tBvqwNmLMjvp9xDPwVo1/MtPTbCGRFuasYV+035h5nyXHCk/jdKGMZtMzH
+saOkG0+IZmzn2Dog/9LqsNQQJ1OMKUbbqGP1PTI+fwvqMkLgD4/J0RYk8lSrBjf5wmBw+X+ks15
gQyDoIyp7XiYLaD7oYlwJghBWEmFToRloX8ItnCf8h44buJcCTFFwcundOd1TcGit8auKVWEsB9e
5ebvJIsEH+uxqlUPw4MXEsQZyi0g3lUk6vaAMMOc5rQkV/R98QtsIYZeqnfQ1S8B8+7XliqxyOJ0
4ONQpGbuVGtlpS+IDNaQp+CkTYy1wb0PEyBLHBggEMEZ1O4FiEb8Yb2ltkFGHPpr6rv58BAE1l6s
uHMOPo1Rk5UdHskouOJL6s8PF49nyhkmgQ9zCE1pE2IRiU0jfauMhfazbQHdjMhus+az1yDJAtwD
BU0lq6+WUbmK10kRFK6C9y5anj0cF+mfVrnwU0JznVD8gBCtJur7Ilo3hWOTSWj0EJC8U37AxAPm
Lvw/a4LvnaZXG7ZsaehSQ8wx6nqRORMuEYUnR212Mi0hGpRYcaAicGBnUd6CXRHrF49UmJdWdfGe
pliUbDVr99jt2PGoLNMGPolHY6CbEIWKzyqqCKoTOpy7oFwyXpt9uMhpITk/7RRMr0ZQswE6HhBY
jArPHqoXLOeEt43LAKlKNh2bcWQ+/o7PARaQLULA7bAM/0udAp+sqvYqwLzIO6tLr/HrmhBUeZ+k
SXO8/NT7V9E2vKar1JL2qi1xuV4Y1U9kfW1K3KLFgiDSztU4Hf4bZQMs9vSQ5o/lvSoWH6EnGm+N
pNkKh1+ZTEFMCjhtdLOrKZ297vD1YgLiQ6If+WlhSifD2PETRcGnSCvfsH2ki/cgSUc3sU4a7SR1
QATPDPJpwAkF5SQgVcNlCt3Od/cqVY8RdA5Hy2AYmWNkjM+ieHO3/8MZvARCfSSRFT2uR29HxrJV
ReCmOFm01mWed7I6bBw5mVinbcUbjRBUy0u5thX6q14yUVLA0rn5q5lLW6g+WWHOnmhh829E0P4P
azO+FEwILfVLA4aL/NTFQ0NFHoVjLwkvya1f3EsBz/6zlaQx+lLTS9Z7AYJg/amZfdv6rguEsCLG
C3q6CT2tnvtrIp+CMfi9+p/Fi4sjaPtDg9CpmdXI4/mSBcXIMhHFOFXPc/Yl0PIu9106qHaeEQ9A
7zQ4CLTsqs9/mNnbYPtOfeQQZa8/3NM1DFHEqBNdPL3FNxrbQxRiegPsiOGVKMN/E/HnEJ8JJxXh
H5H4SY9Nj6ySe4vEvCcBb3L5wSI6PNAWPGX7sRH6gh+6eQKXK9zTb7MQJWUR2V6vR9auYzcYMbjn
gemDEuIBGx1WjKubZuL4Cdmtwr7U5b+OZZcCg27X5FwiG4WdxJqNES2K6F8wWgyRby/Wfh32sBQZ
TF688719jEw1AA9kcZ6+Ot4b0pBveAI3OwoiKEZcuxdPfPVYVYbC+XiqdwtQPzr8qSXXTJ8JRgI5
cRTR6A4R2oAHmc+IvuU4BIrfTzh0FhORehADHW2WL8ngUhETokpH0fPiFJo9oGrkY5CdffDQYNdD
Y3C5QvNjelFHA5XwgnL1XCwZaDZJIO43NNRnA8mjsw8wZj/A2ae73htJDES6rOTYIxQmQs196W0w
lQ+69y+QTOLfcm4B3Z9LsXWP6jcJiau8TssVCFHeKjYIFrFQkkApw0m2YujuOjR9/Wm7EUtgSYsm
yDqbHRssS58gokF85Kh2Fm+8yd5Xi/JGsdKf55aEBzppte8YZ17ai11o3GmLPHpNNfkXC+t3myz1
eMkOpk+X8u0ulHqeKgddWnp+/K/kDNiEO9Brm7hXMTIIx/1XDLcgC3Uq9OnMfE91i0vK1HdIhTi+
IszcsWc2YsMTdwv6IQyKOQ4fQZRXmb2B64c4QDEwuFPM/oZMXQNuAwrgP64pWWXVm2qH/rSVizXN
lk5UDAbdCmljLFF799W8B32Salqi6fnjTD6/YxJ+6Ds/y9wJy+JoqiIu/WA0EqD3FpsMGHa97kz+
2uHgUWak1Z3jc0ZR0cB19VNPGRu7E1I4F65pNIWL//Q81jGmL/n1gJHkZnaSNuR60GFX2dJbGHNX
7d3zrKXcKu4/GL5a4+w0WEAkF3tW6BKiSZB13zFohZqeLzJjjW9sxeAlpmLVmsZaftlKA838EWW6
YdyB7u6yGC84+F6S472V+vsGUZTwRgy2PynBxpm3jb3X5XeicuKO2JesBH/mifCyxcAbqhOY5vYv
V6PfRbp7U0S4e2T2/rGQUOVVMw+sHnXnJtlu+/P4XxHnVKFta+M87v0dJb2IfUVCGJPqn6kPzysO
2F69hg5oIeUWtpX5PKzAOHorgbRYOzmAkbVdHkjPV9IKN3AUJ6lwy9upfhr+P6UtaTeA/gGJnYtm
fxVRxt4boAjwPpOI/Godyo7xlDs8wZ0BdJFJejwYdNYBR+xhJZhiTE1Tdwa0KoCeXigfR5zxOmjL
JECp+PQxLWXPVLVIPGG2wMS8ntjCA2so2lp5eARQOAsoPgDzuZ9bPyWohhqMjnVomOZGCKdTM3aM
gGg2XGKjTIOAPb5e64Yao8l9jY0q8dbSnencjOXnQaVN0H9Tb8IDrsRikrPQMseAPxHGVj77wAOP
tX3qxY97jOZcu4w3YNngpIfRUDH4GMTOt69hAZ3NkjZufLRnmB+FQv4QEH1p1IA4llsLZjnKZalx
UuHoxSCD6xQWOL3D3PRbAiN63VeHXWdkspdqUoM0Uk60C4UNMVRiRTbiwbOfdSjUC+wwiUoDyDj1
ynrEeaMh8cifHgvQVJmlK7TC29dvHnvKnt4z2SpOoz4mjeO2kQRFf+Fuy56uCidXyJqNp5NdmJUx
lZ5Uqydrf+awBfcvcM6q7blQTmdS6Dmw0Lr3zpvx/2rLA+3hPE2ZhHu2WTmy5I9uwVTgDW931gbv
MJSTCRAZU3qKpafLV81aAYdiWLIOtkzV5O02vcb+lnsnE3lyFTdkfLJoz8Upzb7BKUtMENDusinc
WA43GZbSWFZ7Adf2I5bcv9i3AMq+eEmkVw1NGRrXuBpwmXiqPJBz+4oGYYJVkrRQLIH3VcaFrd24
zbtOPEKdEDOljSHpXXDuz+kxpF58DT7YMNsyQRFhkc+VZeeW55nDMAP4gToJKSTXXI0U/MweoPz3
IQ/O0+kY/zYI78hTufbrqXEQvv2+jQbCLGvstxPDqE3SToRMG6yIKKo14R+wCoWBaTOJeSeovtO6
CdCgT+Svp8abiqsMDqAGGXWlIthpXW57bj3YcEuQxZ8oXA2pbqQj6qQU3sJEVERe2aVDqAh0Ua2g
kfTfBi6cH975FF4+qC/P9R/kRBsp/Zf7/PgAY6WBPQ449GxDqoK5p/AB5J6ITQs3QSf7L0emSNTE
EMqPxe/6HpG5hvLjAwPq4AHbvcOIQ8hmLHvy5I1qRz9Siz3ppBmxCsB006oavWs4c1k8G31D8eB/
fb5VkFXF6BrbR596gUMVw6qcltN3a9pSLri81sJN/i7+qV/p0yUyXPyu2eoTAJkQD6UVhPkZlQyd
E0uaw4hiXqPM3Genfr8W6a6wlV8ogSyIGT1Jt7jbXUgbQsIrqyAQVysiFEipO75lM7l/CzWeEqoy
x6Vxn/YLdSW3EQF2XkWBxyHQWaRCac8iRdd8LR/Oe2dYaCvLZprtpRWIvaoq6SVLaRfWRrd3ahNG
HCdrNcmFGQQvpx4u/6WIt46Tn/m5f/BvG8vwkm4k6lnZHEZAohTphNs0vXXpB7hGRecj7A1Jo98k
Mom3LItWARMH4Br5WiSxpz3k1iiLUDppQUHGgBZpWxt0lhkMqUOpAKZV28poA7u5keIGB7dusAjx
LvfTWGW+zfrMnIxDG+wdWdklTqBKA6YcyVSaOz5qss9BvT4LRFUNv5xVpqPmvA53gVjGastyIrvH
+5sZEkcT9Y47o+2TI9B/1P/Rl/sV7FeLiLlpgZsrYOplHKhS2siFKnkKipu8EWPN+lJtTdu8+EDY
jJlqlpyn9gRZC/QSQRunhAZqhsuNtCeaaW1YjPdlCYZy4dTpORtMHq7D8Eem3hyH/usyxM+1oRiN
8px6mLAe0VDlIs1BF8D0XtnQIO8u1gHtlaCvBfndhWKe4RkM/M4H1K70YOgsnWQrTvr8LS3DDOWR
OuKZujJ2bcD0asIbdeVY4k2dA2lGB6ohotUmB+jkcvtw4ecnVUlC4A8/g5nq8Qkl9FrmbThiUTPz
aBNBUNkXghQZr/rWlAbW5qfFgtmw8On1kOL7GqmvxELYAcAPhjsPnZoVT85kynnCSK20Wr09ZVgn
JlNkG2cinrBpXP5QmmJh/nQ1DMmhX4trYVXAbGPra8l9UkxEmX67pLYbSRErYCgb72SfdIWqEDLT
F2jUJgi4WHqab2w9WVyqSZuJaCPDg9Vre/zf//PLvoEqonQAEELrHLYBpFu1AIwnYe8cn4MFCLzO
K/nJbIqfTGI4iJSpUV0J5kS5vOF4t4BshTuK1up7gQ4XEcaflCVaeaAh6nv2cGMkb/fV2yXVYK/O
GMAuEWj097idYVWwvoRpk/7GLf/I9UA5XpVgeiCMJrxoTD7lYDf3VkJnuPT6SR2w3yB3U/06amcu
6nIzEHAgzKoh90cHn7FQk7mAndY9HhIEvX2CgXZF9NuSHKsf0XWb/B4UD1Qooc5m54XzB3BazVZX
/cTeHsPIfaSkeYz5x1vbmmKpxC9H5M9soOQxiB05Yj5HpS/x7qMUbrnbISn05ZctWaRuZKBZN3gc
ERLpOWVIhHVqvdlewOa90U965LEaJI3xY/2zBu3A5AjufUNXsY7eJTFhpanrvB/wZxBXfhFOPiMP
6vgmr2k4QVvFckWbyY2GRrFDnlbxWkIepaiJYwQlDIn1M3mZfPuG0mzoFpW9jfwWLhValRq2+nsG
IWEPIfx+50VNZEYU59lsK71a24ZP2eu9TXv2O5Zhtdb69puz60gyRLmFcVlJNPaQj4KQmHMZJ9SA
pEffVY7rO8S7HzN78r8+80d4UzN8+2bC2K0aYS4R3pL7Wulg+8OiEa7jp2W+zXQCkQE+/7EDooxu
J59ojrb19uAxovD3ECdIwpo6geNUH0J2XuWLemwxQkeJnvd/rZjNtkqy8uprIUYCo8uqs+U+ykEY
3x7kZBUc0hKDWTsMxT6DMickdbmcqAl+H6PDJcq2t5ZJ6X92xkyqMPEPWLvJ7IcSiykBpzfn79ON
76dyEC3ws8FnVTi7UKsnYNEY1I9lJwNaZEo6HFTNiNTFXw689T9LHKiK6qtwDsX+KH3QFemZjnhC
P+VScE6dWYdXSDDYtaDG2y2fY/kuGhKiVcG088ga7nQcjGNcDfAIUJ8SUxUDSYwnC43lkCArAzSR
UGFzBKRLPq2f4aUNQxbn7geMthKunk8dQ3vw6cIxyes4ysFXLYT6KwOwSVjhGGc74DMYcS5Gqmgd
H7MKTnJy1VH5/0l6ne/siwvLb4cXy8i7LB/aUqb6aD0Dk9hsFK3GqRR662TW0QUCOj8sdaq0HUVd
R6Ut7X4aaEz+vF1ivpooUtHBGdiimRMdVLXR+kHOjX5RKCVYz5lhLLiWZWp4cRs10ChRPSE5PAWE
v+zi262KqDS3fWxquXN/9AA0fOkN3z8zHYGvBw73ckUtyf5g1j0DJWfNN+OBwtgtSOCGv/33OaCx
avt2dl6OS8LpNsqY5JrWGBkDpNFtZbyMBh0li2CrOjmec50jugPFYhVpjYTt9t91XyYTG96jpmjm
1CccawVAGgXlcNsjOfo++7FnJD5uI0Ih8NRAh4Xwo46RG9l8OJSevlvkd0ZL7XEncBIEKUTCZr5J
brbrWRejfp6IBKHGbrkcfML03CUmJvNRtYE8j+JiUlmSex4UrAlzQE7wDP4h5dqLmQIEziH5VIb/
wW88v+ZCUQP5W5ev1LN0Of3BB145TuwIYObeN0HgBaEBHD5hhIyNopLcZ5Y5X3ZOpVkD8HrRv+dO
L2eD8xKiYp7a9tLOQ13mnU5eW9FTrXZVOPz6hFROXTaVcJPdqo4d5X0IY8QHNpBSUi3GVqOGiBKA
Y4YSrkhAc8XY/EDAuuse/pR7vPjbU6hwzZMt/YE/l4rbBZaGR/X30bw4pVr9M2EPZo1TgrZsr710
m36DHuAHCPKZBAQylyfp9GbwG2LhtwVSPtabVAUnqTay6s1ZRwXKxORMluYVrokV8CK01tYcJxgb
0cjJn21C9io5+UyZ+40UGT2HPIC0e/ysxQMl15+upB+3NneImV8RG8Hr6BRT7t7Mvld3EaPneiJc
QlGBczuKaqitmfqthn+Zc+3oss5m3giEH9Fe1fWk5kUiwbB1rsON7gnI8PtoQGnfIZIY4S+aHxPu
OXHvcjUd7fDA+Cz75gBoF2YpXN1EruaUtGcPQnDS3ApB1XecSaH4izrCFixZFVy8qf/Lj64sb/Rq
zOPO6JFb3un64rMI3bRQdK6QaKwzHdesw9Bq38AFj4jAh7Vb0SYsJnWMgqXSt2wSGE8f8RTrqPeu
/PmGRRQ+BBOSMrkSoT8y+kYQ0M91i9qsW0wRlu7XxF7FxbuB5JJhiNbdvQiweST1rBTnDvnNE1I7
GIHvOTc1Mnx4PP7ZXn2b83KdVdRK/PZkr8TGqqCdBTfwgKk9YPBnws5pDEs6bZvOU0YohGb57R6n
mHyUJ6uD8c2maZgZ21pkw/EVir663mQYdXNJ2vJiyjXeRDOIgvKZJgT1CZmwqjGQpPNPm6Hc9aqZ
vrehbxeUg7JQDXdh1/fVd+Q7gt+NEslwoOMHVVU9YRvwe2N3/my9eYwwRADrX97gziQJk9re4PVh
t8l4eEsiY2F69ZYwGwGkvxZx1JYXcAp9dPWuTuFXMtqTyBOje6gLk0BmcDfHqgk3JXpRPjZJ5gLF
fG27ciRA8y0w1MFtb0Xmjdvn8UcM2ivYpsNxfMxTQvS+s43slhnkkOROW86IULeczP+Nhcr91Lwh
LvFwKuR6tQ/vFFCFqXmMVkTcA6KOFqebWn6b9uKMxzp8UVyh+HS/8Ms/iVsbGKBtXWTHoRkaUtDo
dc1fc6KUzTszRBD/2B70noXfZYx99PZRMWsB+KMT706SGuCn0E/x7n+ynhDPNFrFNsE83vWYzpow
lfbomQhksKAEEGf1HKyhEa4FXTT5k2VRMe7YlhaApirPyzHjgPS9rZGB7Zz6PBHXowxGYn8xsY2g
S6KVObE8vWnoOeXQGj3hySZ4tCVSxZ+EVRy6F7e1eiECThaJhFZWApvTUjUBcElFjoS7TvcnD4da
TaA2wjXB7fiobmwuzrgmE2kEgFt505jf0Sv9Uo+ogJwZjmNg6ZPqaJQta91azWFxPhAO/dlGRvCP
AKu32UY2vF0EK9LVDkagNTdgdlXkVi9EDQKxfzlZwtfDuDwIt4deTb5u1DxiH+Xy1CG1SkWjmaj8
J9qKI1jyYr+sI1NjQiyOC70v+QaE/FIr3JXwgB9dyjxEcsvt/1UZJNzX2kNq9YqdTBWdFzFi5wQu
l/McjheU+gcfTkNjPrhwGS+SmmlUGl1gklGRt1mBHjh1DMAXjYcCx9f8uUsKXjD+UnFbNikHMcgG
b1ebGR8gR2s+R8ugNWAtB2fBtHjjDSVuvKY8KlBfJexnpv+vNmcBX/xiZn98af0SUpdFDuYWJoMK
Z15m2rr9zILg552TaO9q7t87WlMZtSE1F+sWckTuRAsYrlkHCWdX1U1Zg/laMa+I+298MVULIkLZ
6s96k018EokC7wZ8puo3exZ0IPcgo75lDp60f6sTvriqyp6dAx6yGTWCJg7KDtKzqU+cbCie3t7C
EQoNm4QqqzBND4zFNoPQc70+Al2yWA6jPZzgWFwJqYqFpVVbFG3uV+UaglCorKQPwM895KAoH8zC
Qy6nIa+HyRURsWc+f1skYtuarZO9Igy5MyAJ1XIF4SpmSDgIwQtADbZ+DmW9iVA8JfCJYaEmQVVQ
4cytnw/ni5YHEngwpAGFpbyxZiwuJVGS+F/ZCYUATYsZSRbfKdqonMU9b0VqqSckpHdkDFY5naK/
AAwGNek8VrDrPYavhWSCDB7f0984cYCDOdqSZrIRZlRClGV6kkUHbp+bHKWVEKeTtaNqSTdinVrK
/k4HDEsVHErVUIJ87cINxkio8F9xihuXi0cZAas34tnpInL7OGQw8RmdB5Ljt5Sz32af1VTXx/Tq
haYOI0AEvBVkbAwMlKBuZel8BUpbxZ9oxBdQbbeFhO8WIgBLnBTj2RE79B+t7QCEPvHXGB6AL+he
zYpm1eTkzRdEhcf5HNbCLp+UBh+PmuoeTPYbSrKD8ZfIUxwGIvv4S7tB8VvZ5749o2gdzRnymhGV
TpkxoCWuY7ObYXJ8mvsg1euH6l/Xls3EEqImDjNN6yI1uZM7/4V4b0B69VcOvbYE561S5/KbStus
HwnMFxWQWaEe9XbPSYP2mJU986bdaBdjZBSghAwjdb/TGh+3JqKf+Jf0lQXL1es2uczTDwxjrkbx
TvV2gcPlWX7b8lE1Sk+MfbjkqvTGX+or/S8jK9U7vRMnqMFoufO+rlBIYe+7BP4zO70YY1lNUXci
PHdilC3r/bE/s212IkgfTMiSy5BFm4zJXtt2sTmkApu1c+AI+eF8irM0LudDQOKOs4v0XqtTcYyp
AqVSBMazRriR465MQfbFZJkVnsERMeIiizHe/jchHvMZahTNjJnGwULTb0MgKxlX+F4o23uo6LZ/
uxN5pBQ7+//XdRmGVg0Q0BjyLjXcrSilF2evKqkP1/8gfWEJ2rBK/YaGthhaRb1jkEN4vrPRznQn
TN4Iwe2TcK4+g6km5gxlLPENXh6C1PzsbWM9mQ6hrVdDpvAPF0JXPqeDQEPuDHFRMVRIKEFLaNFe
obHBjcrsOcbNq6viLQL22dZxfz2akuspXCjo82H5sX/9XMSFWPmM612Gw+3yWRAMZXGjrPt3mVP+
uyxlUm0VSJIjKzAA/FduEzB1uKS7sHW0983bfa48Cf7cduWKaKEZGfi3kNcOJCZ1KOOuZ9pmDDL9
kgQG+U0N8ld22nc5FyTr44bSunz/01lDDTN+B5OcKeUgh/0ZeX7tbW5LxQ6+6hA1X9lJPHw03RI9
qWZIyuWKJsS53+FMsWYygmn3FfPOAwxWulcq68XuQ0kfbf6G7Cah5/clMvYuFsch3DaJqnQyw9rG
kdg2PQIul4LpreAs9OtFYGfUY4bEXYV6zsgiNawYnUw+emPL9+dfSEfspE/WdEPkUkT1OygO7pHF
V7igRBmYy5DZDdnTIK2UnI+uqNEOHkn8HcKJW5OszmQybvS5ByaFEBkzi17s+Ax0sEUdft1JuKoa
xrd7Z6P0WLyD+mrQGIPD9tSpHBD4EY76GhKjxWV78Ah6N3EH+SIlcmDQN8geth06Lg0thERAqBeZ
h/a2JFhFIEbilNzvMSA/NW0ebuy/EhpLx6/77pm65yO0+usUq3ftzvreQYADaGxiu7YLLq+69kkC
n3BBTrxT3yeQ5FlBGfNhkXTnawHItey0QJD8Oq1SxvxuksQ06NLdz4IlH2m5ZQG+m19JPo5t4fBS
qeN58GQm4UGr4bMdPPqsGKbhODo1l8so0C7htTK1b+XooRkVZ84h0FwYJHCUBY9BUmUMt41NSULm
U+SicjUZokwFpNECzcLvjg1QrFN2dtu+HRq0ov0J3EWROXLp6x29rfd6gOhjunzc7lxgB/2xBaDf
PE1R4VHuRJgKNrluTFSOgpqEdgce0ss8xTKXsTM8MimjDPLDnWfaV+ByfQexs5FYutVTofXS7oDe
hMKYBLQzOFwBFt3JRo/XdgvDnnFpAyClCD8UU270bb+/aBl/txEQrDw1HvFpDHn3omKLB50YHBi3
CFa2NDCB6Cmm9eEL1USpAI4OsG95uFE9NzW2jZSzrDw5aklttLmOaX0zoflwA1cr37p1wnNjuziW
7DpEVOwRWgMI/isZfSwM0L/EAHo8qg/fmcrg9o44UfJZ9KC4zY+K07pUDNd1j55THZDSibgBzci3
jgpupb0l60iCn3308WZ+A9sK33cG2SsXwPP9Numih8WjfjCUhL0QLG2/GPYfgt4lmlxPzH3qB7ym
kApDTqERmVAr5nyBFwetwutnMu0hOJf2qZUoHinHcLNlFECnGbUzJrIkgOXYfhfyS3rwn7JoZGdj
hcz7RXoFzazNg91G9z8Rk30ASxBbIJk7rEoEKfQZaqEKF4BqUvc/xXvTS3PvriwV/bxZnN9qj19T
JR6wR3fglL+908SrIsgmdXKXfq1SMoIepBX6G7ZfWEpQhS35ybd8xJRvHLQ7CklMf2658JMx3SNb
79y6ZMUSjwgJK+RpgiP42lFOMqInkPzTFvdzBF34VTWxIyvSrf/aoKljgAcC3hyxiIZSdWShJv4O
T4vZXcdiT8/wg/zHkn6A0J+wkKFWK5XFZJF3kKe5sQp1NXSiarrLmudG7AeYsStsZdblkFlMprwT
QL38LkYFMTFeiHx8EsddTRvYn9dmePR2YnlZZMLCozpJ7lG0OhECjGLBMb+A2aQ/1haGv1tvMdy2
cMO5leDpWP8D8tbspa92m3HsPFMelo1aCRZdkBdlLrLetQlR4Bn1m+7DJg1nskUBvcNXdk+eTDCk
zeUR98qrT0O0U9r5UmQo2Js35Xj8O9HFX7ykre4YOB4/4gXiQMggy7egFxdtfZL5C1SFIyW33She
FOUVT2XmZt4U8u1cf5+dMBDsXfNr3p2SpSMrxuReEFkhRs/1PPv9uGnMlrWcQwD1PQ3Exwx8btH6
pa/DkE81qLd8LapJInlipIt9TgvADCUkM0v9O16g/p3/eRC3yVaJBS8YMM2fCE53FM6yj+uQvtdg
/hF7ZIE2vWX2CVS2loQ/Y9BLeckGoCp5la7yujNpA+sH99hEDZ7r1A2v6ZHtAtSXDQSpIC7Rap4D
ySGqOosecgH76gJc8pdexeJY8WNl3NZxtHtAaIJpdiGlIWFWOEyIzM7atYu+MtqkgyBkhZf5vLy6
+FrRgemVChBsqB/X1gyYZ99yaxI3v9LYvqGmYnN43BrFGrP+V6SK1GXT3MgILqb0BY54QEYdr52s
cGa9peqIa5l8dMc+WKg4JUAZ9V92EegHDHe3oTUdKOZPSbHYInzrN8QBYJaWIz2tEPntyQEP4Dbn
Zsfbd6nK5h4dlFU+MZN4VUCUsF+uALIdtHr1tMwN9kFZQDn1zwHmUJp8rCPVvCVxgzZuH+Cv2tZh
EUDby/h+ATnXRA0KQx1pFEAhgROwmpQQUqveCAqg48EY6NoIZjULsmiudB4sMqe2x74tWzFswFsi
qTR9+gOD7q5E7pcR4gYjAtaheE3gkh1iCwSI1cid1yPLVfgMihLk+E/C8cadww72548K7Yy9Tw4s
3qr3AUdG2jHq9WbziX2+7XTyHOL7p4IZsocuoU9AO3bfg9plvYW5RIZd1Vu9m9IpVMgIYfTLN/O/
3oC7rIls96uRHZ6LYtPfPCNSTZMMsNCf3v+s9tLDDwcwqUx0mOSzRE2Dh0d5CAxCXw75xDzbCwg9
semU9xOI4VdtcF69zfMp9HZH6C59yY4KWtfgL9WHoXrCYXDXSvM1ooVVNrYA5NcADK0bRnwCTuyK
ckj5GMxjj+/WyYlfBz1bqwag1Mp4cxCjx/bQEO9erBUHJAtxls6YEVVNhPd60sKCiPqxjtNmTz2x
kbIVMT8XJTyTUNpLdwV2gUhwZjyB2xgPb6FsKsXO1Xatz75+DmAvo2mz7yTwrl+U+FkUqOHNco9Y
CXk8mw4RvSmuEqkYF7GDyO8Z5cfS4/Wukkc8N6QNqAf6mG6SVLRSvnuJUyglgTg7jPl2F1+qGcbU
eYgVuHdiBVERQlCZ+NrPd1GIBe9ruN6hS8v4HFu3zQD+32/94p7D+wZhbTyESi+iXa5o92KAVSC6
wmuyxiVXmOVDog0E6Q+RM/a5yQ7Abxe3B/R0WpojpReFjXGLqwQV1pQsaA30vta+7Mn7hnQtxcB7
C0EfUPMLExGAeT1S0wr44eJRQY/+BNC31S7f8+HOAuDnG6NMGQX+dDwtMNR5ocpbG8WoNHScRaPV
OLKzXS2SRM77lPLckvl6YYXn5VBHr61uSChxDV9auSDg9QeZ/KDGCURr4Zi8g+DSnIjyRZf7AyKO
dqhljNbgN9pZXPZ6miHNWv3itmaqmlg3g4NJEMO2pQMBfDyqb1kgPvMnqqxv+XVxAZArpioYY8+d
rMqvUCv1hXu+t8jMOadgh5e2L9xQjN3lQVmIJ2zV11HiBn/J+FXSDtnpnlFFjRuLnOjWGvo7+SmS
4kXMJyD6kfv2cfdNCr7rZPQ98AIHpbBo/k77BmE/dFUP3BP0H1pS+L21Ch09kILu5WvAlkbQ/Da2
4Q8FGDsi++LHJZsaxGwhVKeQo/qOXyS6zW7++3Q0FjKrOmL7BzCh8xt/3gJVxslB6LHevy2fc18y
Zpwi1llO/BRulcYtODkRCOsCFIRqhFgPGRB+JrdhYjokt3JXoknQFaediy/4tAGwEnZJqqXQhk1r
kQZMcG9U6qIyQHBZK3kYSqFUDQSizdwR4uK0t1ltg0sIG3aBGhcgvImaX91GHAVeND/wN/B4FSVI
DsR7gXsht2oYmuIqMa1YsTSUVHCuHvqzh9VuQrgj6ELXWaXIgVerqpoVept2Qi6DrIcD89Rj913/
cAdrhQ34uAt9GlAZ+rKRJdwDeaXFrD53Jx0BMRS86xbfmMqeZiixcc2L+nb+X/t7vqzDfAg9DH0A
mkoneLXI36OSADvtidpuvH+B3OrsVLF8n/LtTn3URaMPMRpEOkrxRSXYI1pwZZ70usjO+KeYDmFv
iTvqMDWn2s0Fbuzu/0c/9DD0KtAB1lFG1/FCO2xAKsvs0vgy15fTNzKTPSHi0nsFpnA7wZ3vhEgQ
qVWsAoMvWpAXVbDGoyDuE6gP7wKA9Mc2pdZaVRg4UnUBmjX9TwgaSvd62OmVR0hucGhOyXGbxNfG
4ymPYdJ7wz9VPOWPE/GTO3qNuds2k0D5IetWpUp1EIljcwNN9FvgPsiKClpc1wm1gslkERxwsfDS
/HTaiHGBl1oFqDEaMQxC3JWHAyIZKLBCfIh9mhMKVQw+6hWwZs/0OFObcqAwW7RDt/hdXIhKcd+v
8ZnRruxM611tj/Rd+Dc2ZREQrGNJu964QRb0FVUcx/VbFLAN52q6fcu7hbNH4kxFcgUju55qouXo
H2VDO/dulkXSaPCNSeY6n9x+FNG6DWrNKRC9h0yVOVaoqWEcX4Isk8RESJtN3hi1L1beJ/Ieauct
bjOVDEudSnpia6uZzAqb6JFUIORfl4rMLqyx9w1pczitAG4AUVdhjXKZkIqCiBXiV1gBD0mzd9Go
Weeq5z/0OjjxRo5PxoBWxfRWXpdTWfVeY1lasVlMMNIfjjIrgUi01+MLR190ytoW0z359WiJClih
s59Qsei5CfnSZAybwQXu/igYHs3VD1rub2f+kqoCgoHzf9H6zWG7FdHleU5zLAn3thSsQSqGaBnc
ZR0odxooJn9p6oTGRcKtlPmywnC8ZQHTM8LTxw5cJrpFAX0rzL/knN/hC7iNOC7Y5JQTXFv6KJxt
daOlgLMvR5pjzg7HuJ91nCanaLZVKiBLUgHd6owQkHhoeReli2kvDBSL/H1MbtyGaARr/Z9GS7IW
asUjY1QfHrNgyJ7aQEtivVLusJznvg9pl3rMLVDGn+CxZZbBLdGkMMVyVfaSkcjnbV+4Rpgpp0ct
MhRIUvxt8bEIAv5IECv0dVEMjuE7S9jnrs4ZvkhrPBuS12QExSvpIg5R+Net2edX0xPxCVwHCImO
if8xUxKANmWNnvSoOUVRhAyksI/6wVgJCfh9biPJBtD1bZPS1uxYDJ/QawVMd7Psz7yocg+ZWUu/
EbyOMrgIpiFTL+gCo5Qr3UZedNZIkuoEwGTOeMwEC7DbaORVuPH3gpUPRam3wsmA8O/U9VxujaWo
EB9+b3dzpFOzEqJivhO6IMbB7zeNXMuzXiwNj8fzDHbqMCYgUd2SlDVQJq8FWcoIMpoQ5shUm0d8
uc0gSAIta7TBt5Rb0Q42WtuRbZmNkPyLuoTz7cOB1f7FmUXTK4v/OFmT0VyExY0MqS2979DwQ6Uh
336E1teMtuG3CrsJVE2dOEQ4Y3jWWn/wyi6FG5ZNA4efYY0x/nCZrVL/+q7dovoz6cKk53moXZKe
dTl73VQORfnc4r4L1AFcemzQToKKWYCTCkEAZ050cEAlLDCjd5oTuGVQaVOkfW0r/RpL0/f+38VQ
BFVqKbZeJG0Phz90Xtk62ruz0yaV8Qeep6QQjOvxtLZQPyq5vWMPw7A9dyB6GTXjKTIoedPQ9zHf
gvthufZp+WMm3l1MAglW7NP/tGxEryz7yCow24wDXDNRLp4QzQaT8N5lrFLqgJ06mYqQH59Hcnmi
HNVopn4hdYEtrj1H77ccnpWPpjJD+cHYBs/e0CoHFbwFSbnEHgvC5k59nvDJwHRHXHEyEgFRDV7p
mKoI+cWXZbwV5V62y4NTPlqaCO5Gh1L/RQUSxYjipZFyoimz2Znr0owdrOo5Q7QBMJFZa/JDjLgO
My9frW530SIFO402HoO8y4guznMsrOD25LafLKYvPvtJnPjDiZEcDv3N7gmuOmGzKyhVSyMig0qo
hmZ0r2PumjXxvaNinunuicRG7NcKBP0wIrg7aJwDvT+fS7GVb9EIT2wWrDzhh5Ge0nJda/XIELKT
OzK7QkUc8Ay4zRWwNeV7u3jNMAxx7PmLQD0MGno9/IUhmdYdf3HMCPFFKrqjTuasW8RVwDLC7Wvg
3tYsmobKpFVIyLaaRzpSHJbn/yspwlWlUiGhdU8DD/mMA9eg18rnItkwoWO2ClsbVzVuCtEBaoaB
yLhK0nt3g+uGn+8PPJEqXYEEx5lRCajHf8+Zv/9Qv0ukRDgJy4lHf6mOkhGawejsDOP2iurOhFfy
+mII6skUwZ8z/Sl9RcROIWO8KfQpWZ9XwIKR/Z906qSTh1wBWHBa5v9ZsQ0K9OuQEpqdTY6q5D6y
7tiYzFw25TDX+zdFhMuS9iTgJc8XVFH+x0Lyv47p6J9ImgxWTUuM2GbTa6q2MCMgaFL/x32LLfHM
UfRRMhSB7mcwzu7KHuWePmIMyx/TsnkzjFuNLfX7ee/NZuRgggkzqyuFQYMoTKaaUnJ2wmmdcDr3
wbkcean21Axw3KKn+QlvU1ntNrsws09ISxnA31vQVtUqREWv62wE29TupYveZKzdkx5ioaqvoZRQ
7N4XtHdKTfP0R93DSj8yENPYjJUh2KN01LDpO2P2xH1UUyVltbGHLfu/ZZgvjAWsM5De7XBvAPD1
dGZk17Z37a923yxPdM9ii/0XOIy5cdi2oEijeze9z4EthCqS61Ij9CatOADIGo+eYXR3kcxdNnz/
wAtXV4fjpG8yTtELKcm0L5vSWpzP/Z8WI9AVUDrmlzT5R5S/24I/vfzznb4SRfdx8CyDdCG7FGMf
1CASEoAlq4xycercXWwagfVEKV72cbFiwgWaJQ+z5HJs9JlvfhOXXEdtmJoALudKNmFRqUmLV8gq
aaLz4rTzjHItPo2TP6SwDIwskUCy2t3FVffAI3f7jeF08a0idLcOQdOe2FgGeXjblfILwAyRl15L
Qgl1ceSa1o2WFUaC142K3FriuHSFk2O8GJlWsQZF/UIfyyRaD4gqafEaPEAKSlLJRFdA+/Z6bNTy
2mGEVqH+baZL7nhzv0G91kcJ3dRaQWTJIn3xT8jjpmR32xN0+lgx7x8QEFxoQkyVaILwUT/V3RtN
Fdi5FWza3b/Aj94sWlnTV1yIHrTOvhB24y3XRr46uTTiMqUfHqSaGLcEG5rgv6NMV/JBCphAckE8
gCu51VS2RIvtQ2NUk8Mxv4O8y31BaeM4XPOMmLKWnu+W+qkok3oqkFIs1cmy7D307hfysqz4fydS
y8wqTgJRCJ8nK4y7OQ1Q5dzDR3y08cTb4/X0TOFzaiFwnoQN6RuewxY6DyJs/0HI9jX9uiIwDxni
R4VqB/3Su8nixmgRJ1Mci796v+u0y1OfHlF+JEQjIpsdEAJsBxWUjS0IZLwGJkgwkiUIIMxDZHl7
9PZe1LUxNBPpeHuUScIVJ9LhxnBqV4vR7sPqIRaHyhnmxr1gwkPuXulAuc/pka1HEpXCxXby6Phj
wR+27A2BCqDX38LerBxpE88GPCDn1TVywiek68KreryMxb50or3YL3HF2qaW7Ju5L/f9O6blPzlF
7RR8feHEyXu3/0sDM2Gartxnzt2XAC1QAD8MF6e69IBWT1qmyybAfETEYIdVGrSaonGgX6w54rFB
hUl6N6oSZYYOS/tQuqB5cj3CPr8lO5RtuzDXlRHdj+ZVteXjR9G944tBvmT7wSJi2x1REXphIy0P
2pN5iT0Ev4zQzcGVtUSY+tbiM8ZlL1+tgZj7aGSpnKrM4SMoejJ0a4XQA2gAZEHXiJ41nkGF6S9f
sj1E9hbZ+PsmrOpHamV4WPyTgZIAKbM/c2kw3NI0UdvU87rMhmiSIhECz50bjVR42ZXs+mvOYJbc
5tDUt+oKtfpkw1L01Sq7l/y2oCjhqWTb38QVY/whxBxcTo7PPLFO80l6b7Fc9phFYtwr9qpsV2ZC
z/c3HglARd3HviVjVUnM2tDIgYu2Tsl+bMzsVceeCT+H/geXTpfGDprnb3VOUZHffls5lFirQJq8
wlQjgBFREvFUPTDKteeOaa9oz4/icia4Kv5UA7s8JOuYxKihDArcY3Y8TqTBcgxdVBnKdTxboUuC
myi5fDUrZiwP/jQCYxiDH0kiHqWzwTRVrrRfvoJ3jLQ5DdWzfp8sMeTccgfAdMtbFJtPX+SpXUad
Dgq57RhRFgG0mhJERaVBiFZboG5JYcwSfGo/gqeKBuCdzJSSwIzrjECaZOJtYy7PLC5n57B23c5a
KeMXBpkiRZt7OFK9yXLPmTaVB0oR623XKDhzYYNpnEh5bpnI0ReMp2oj1y/WAcF/HzubJWI4z+vY
s8s8iYCe+heBALnofvbu96VrwgtxXOwbrPk6Y6RbLTtGQ8bXarspuaaEu5eOC9dzhIzL+6UYy/GQ
TFOvy+lMvfVYMw8hRjAgaRoEWW2bnbKZPrFAktaKP8nMUUjcukisRtAryyAWuuRrxZWn5zHuTxzQ
jkNxz0nWp5INYuL4XgL9BqWUZn3q8gcyg9lmvS5hs/lAutQ6ZlsS1KcVtSnt9YclkwBjBUov8dsG
7uUJwlXsNwR+KyGBoVJsAQvjiIMlH/a5kYd2hzx3u1Qd1Lli7tINJnhalEFjSP1HOVh5ERTIaCLh
Jlo4NitaD2Yqzn4I34b3YAQOJ/DRR5uaY/0o/Vg0w9GNjd41s9TEZEXIO/fV6COZyTf99fUVTnNm
ANO/FSBrt0H4F7mfsoW3CIlXYmpOwuTqXCSBL9v1Yg03XT+jX1WsDuC2JOVgdNTcqOssXSERmooi
M4GNMucayer3rFsIGOkjZd0vrVlOfbk1/nA/GB8bJr4sHm+Bele1jH8s1HFuR68ka64Uiqk86hL/
nNjZ021RwM+wXvUxEmAIP6VQGV8psE/3bhNDdWQixcrz7HfNgdlgGsltMLiKpPhXjyeivRkG2NBi
Do28P+rV3R5k+osfBdta/whi/5PMbkhi/klfyUQvNpKlXd7U/R4J5Onrc+ttxXl7R9jYKEReExuz
+UXjXcsL7jKcWqAZUBeaKbjvlVaYCSoluCOWKeLtBYzqHS8SPNb5JvB3AtDPbyNi8fs9kgw+DiZg
FjzfjsDOdMwwZ2LtjUGkrb9/W4ZP/lguYIfOV1JnnJH0IPnkCrl5NsWkKo8ve6MaNuAOLWxREPt3
9DmQwwXSp4vGBoIQLGOXg/9CMbSLeuiejvyszrRoSxzvKb8oI6ep27S2dHgy0TGOXeOcbTKbC+am
XTGDpxiLyshfLnJfMiYGDuH0RhWoEa9kRCotXq3AmyyinzlLVX/LDupjQCYsITokLnhQSe59VPer
TvRr5zZk3tJYP3uUKxBHbFfnw+rgdGq66MmUmpFE2xqjEgvDFCGGu4p8IIylY4xmYE46Jp7YwZej
/qsWBp4543foVVO5Nml3W8e1H5QvdRNyy0EK/PzfIHIJKYs6mjpVB7yjZgBqYQTVKf7Lkofu+aDD
8KXRYkpaEO0jaUx2RgFBit5gZ5nuUDNlNSWp2RGRVYQ/ri9/eNt/Ax2hUc/BYsF/5OthT+3EKaI5
w5z1m1/krlsceuMDKVbYw5JAdW8wakl4wtz4KoVbfQpMfj3u+fWbmxc0vrzhwtp5qZhFK2z2uIuk
YV+RqXsCnZf2qI/pjz5wT9YLnB0cVGKbHIVRJE81EkbUtjrO2KRQxv+pcPLYLYVDBkpRGoggVYWv
aCBjO4uOZ6zA8e8m7o+7RaHu2vPmqdKDn0AM9EVjJz2qynblemw2RpCZ5s2z8ZLONe42+frlbiRT
+7SfHJxKnJz6UVZWP1lkebnbJvIr2ieDPB5hdqQBKMjH9Jpm8iA1jbfUq/8x2em4+yRbqoRd8WdA
Kgnh/swRH+6RJjFt7FvZAf48V44s/dujLf+8wPIVpf361ZKc5sM4tTUb9mQ94sBS+lqnRp2LmqC1
+47of6UclUBz63V6Ki5QO6atOkRTRgBXVwLXFHgr6V7DLkcb/m7aIoPlVggLpb5xsmhSL5K+2LUs
X5jTsCryFeqlY88/t1AAYrRk0eyy7aEFl7OclanXPBLfE9nPu51WcDpQkS5agsILdnL0MRLkA5Ws
TRxHdILhGbCMPDW7oJxqNZyqVXdyeFVlKmpBsrHcVI2TR5LYI1ll+tHH8R9qUPL7PC6fv0sW9HO+
upQyvNOvJASA1plAMoQt6huhMt4ALnFYHN/gjnGhiGk/SRnN68XnbsxEfjEAN5WUhbcsc0o68s+V
20iyQf2d4CXFr7OxMeFzYQ1eVy+Hrh0AzlBFJIiXWH/w+4DzzIuEVNOutX0ZdfWpS6J6NkRGLZpC
4ClRkSHAUdosOh5/XqaQgI5Qw+A79GRVvMYH+p1j2A85ZJkkwwrYUgNFAUuWDdvgnjWO6P21ofLn
kKeflYV+3p4pTk0LOFgB4DunFW+5xtDTcwqBsC/cr19hZfL7ZEPL5eKfLMxBFc4lJFFVI1F7i8GA
DvwASTeePKvXo6KqHJyYn/YFsvtN4w5ku6RtQeh6ejkde8Yh6oicgt9DLsvjBAN1t04h94sblxoy
asSXql3i5QcBp5PkNKUs2cxOTOIZghsgq8sybDp/QjV+OMH5+lHQxWN+SOAEYmoMM6qFYAVAsCaW
iHMdR5Ro/IWaxRbLd8EBmRU6VCe8M1QPxF2bT6TDDz+KH131o6l558vjYaRrAg0y/LzgpRmwsyXm
NpRA0tcb2qr/nAjIQ8xcv7Jyf1K0t1mOkpgp8bfpOqMOcaDAWRj/k0Slee2ob/mzmU+hnWElC+Ma
M15lgfM0CAn9eICkMTr+taSQzwImF6URnzTi0uxGRjakZxGh1QSRrgdz6GuCD/zzDtgL/BDDRDfH
apMZWIG8J2c6+IPU2GYfYq+WQDzUsQJDxrj95WdHV8t/BJl9SNeywmZ0yKsIzVrlto5fZes6w4x5
O/XQtaWZBVy2826+D0D8S0zaZOemmG/ODm0XItoa5ko2JjYdvQSvcYDP713GP3PxDjqL+CLrI4UA
gxEAjv0BFWQrPCfGBRgZn/nW0/WeSJbQ+ORsr3Qj8QQ9W9ZChB/9FLgOZmb7zaDnc0DhckFWobo9
1pik7FCuNpe+gK0g6oKKigg5hiupbnUNUmU+4S7mkpYtb42GbeTn2D6x2OrTOe+J5OhAlDD1k0XS
FSz0QQp1NpeW6XksE2zckkrS1F1X6U+4QmEhiwBLH+hjaUGMa8rcz4YG9ny8+e+e6xf4rum07Wbb
NiH/cmSF/cM8P6XpLrvYXz0rtRaRdT6GArCd/XNB9tdlUlYNHmxrpRvHdMBsMsMDa40XYIQPyA92
jDDiRQpFv2O6TMDT/sRySgSDQb8Nl6H/ldQuJBohDrlzsD/XUaiDI6mms1AcQUe7hUTd/QrFgY/y
aj65YH3q9Srnl6DKoGs2k/egYHTFi/+uIPVhztiYV+Vza/ztzA0b/K/eG94Ow2vN9cYaxI069UzB
Jqc+Z0zupVSQ5xYoXMeo3so2+Jj+QWiyvj4atSPzyONLWGbA87Lf/dCHJtabrnDBvskyMLKR4Izf
STO24gp81Eooalag0rnfCS4zjLEvJFXnKG4lIVJ8jX+uhZ1s0NnRxyBkmZbRInSP8GSriQ5mBaey
oUU8siKNiHhyFS13EukH5gG2EjZ7vrp9q01jabiOL74GBZkN8Rx0Dn+KQKhYhHptr2q0BlicJIYf
uFZQVFSCjia3NO9G+VlOZg6GkK9rPRE+4pl1EWLF2HWcyMjAWpgw+BKNnfdvroIQikEP2grpwoH3
EQoE/OWm11IWYFjX2SQ5rFE8peIIdb+eJZpWHbZnIeCNZu57RU2jnHpU0qxQZMwDBfHmVUkz6XDW
KSHShFd1ElZ50vq60m84Hc65rNOvGXHjMeO+4ciW5176brdmxo2YYRxHueiRGFxtipaLKzv14IEg
7s5J2Qa/PR+4AiAfNlXPc0JOjrn58rnS534j3TPz3m3x+MbFAWE+g5NmZ6K5HYXOnvjfKifhZk4c
9eCO8nbQpch3YgnrYCglKvRNawIDdUiBFBfvToXs2msebIKaTME26j0mrcCVEaN6RWzZYMByuNrx
nhjarvvoaeK8ATYdaOmOduALkUGfTyRwaEsLX5iwfNhn0oxGyzRI5qKc1LriJMK7SwFbfLVt3lXR
+0GGCTL+GbjKoB819Rm4YUexuqVb7/UYaDC+I+1CN8mHYTbV5a9lPAe3B/icQFkE0uw3JbxdG6cI
BZla5WWPkJgfoo2H6OsAGjxwRgdz7SDmj8wZbduocrJ1LJsh8r7IGR3tynCiGG9is2I9/t9w3/hA
ojuihday6FU0vDBxdntt/vKAEtyf1rh7AQED9ie5ZAyfmSUn8F32/GNkzqxD5rkw8LzNohGAhrD6
Re/4nCI/ifsF/1U84gdgEL4mRUsxDOIK5IkrIFNQvL3HBPmutp1ueF8LNSdxGxkw8cEeCl7QfICA
/Oq+JkAJIGWTkdelKjg7tNzh0No681lxA9iVfXcjcZfOJsOmTn8EIOOWNNzGHbSNVYPagjbEjHSy
LeWr0qOmYcmwePpiKv9pNyKaXTXQ3tG8PFwBLN7qaWE2/7wmfCziu3mgWweEpdmui90p5L0ySMNA
bbb+vaHL3A5GWN6xQ6XppfIJ24lQ1h92grnuwd6zP2zKB1QaejIdluxo3Iheg/rdt7EJM7fKJUng
DslkwiCHXX+EJihqqtls+mJtp2f6W1Qg2qG4fUba+HNpZHuvgy59+TJtU8NbkO1RWz57FEvz86KH
WVDzYcvhytupmNUgwWw0B2YiMlOkLNKhiK09qcsHYbD3FaN6l1w/V/GKv/18EuaWd5CGUW4sw7ip
9kswdZTDCEHoXoiTYGL+c3dN/G9QhP1bloiamATTbIpeFG/X7EJ1ILXgfqG+b1y0nNMN+RZJBgNv
V5m8VPph1RbWR0C6waoHe7d0Q7/jlEtdJCfMt01jYn4L1KT8PuFVZNNT4pAxi2KpUQH5RqHJ6OX3
aDQB+fZXJ1ID4uCvz3Ta5XikN7C4LCWiHMUGCXU5rOS4yjmPp43h1Qgntu8DQJFBA0hL3PGae30j
QkJXEGGQs7QoplAnyPb+sR7z+7iER6j56VjaSjBX+GkOcEgdkJJorWPynJqa6IbTkRLKClvYyANw
vaWiUzLSSCumbH48stXLhDxslMS7+HKspKUdUtVV10ZC9gB5iPy0xwYmz6rAVqKUsEmzTLdFGoTt
rFvwrYDupvzmlTPrVUKGcc1rsxSGOW+G00d6GgBWY9S5k/OlqaNeAxTSYtG0pkXnW+N5Xwq7Ci3l
fHxzwqOzjRQv5meHZglUqWX2gQNzEXKlgrnqsZ4uGzkjjQ9K40VyfgKNn5xLWLpXVZ6BJTX9s7Y6
fVClXZ0GwRiG/lOaguUyBa18aHCr6+2hFrVkUYOudIdXBBu/b7o/n335yh511+LY6Z3vxu9znnGR
707mtN6WkBMeUyml1x1/1IUXgI7vkGXWrYXGAsGv9Q9rqWWDg7zQoKofi8Ix2rZ6hcHwEBPSJSv9
2RiJhW0OKNSc+1PcUWitOsfxJlypQIdLNoSA9lYhQcN5z9jlfffp3eb2P1VztIvN0pE2etzyPorV
FYhE538v5xkRqQsW+i5agIFTnMEa5ZzLoppnkkwbI6sx1+IdSG8mFZNhot9trCJjsYyCQM4W6Y2H
A4mmmWm5IDjNsDvIb0ZZK5ZVOwNIGKD/w/lKIbLWeMK16htnV8clmXsuFtx7CgjJqv6xWGnhH8hh
+oTSzZSaePYdlHdqR9JQUkbxpmySgXrytkZLADqvMRr9MtsbBRtoW+7QwY+RuQ+zq3gxm1pu9aDW
5hg+PytyL94TEiUMrIa6dX0Ocpkr4glghLPJYjrFQcHUv+tzhJHQZeksXY7Mc4ZegpBSpQWJv21e
D9F0i0m7fsBgTflpvnGcrJTBP5EbQTqsSY7N1yM0oK62ElwK7ICL3rt5mtPvPhD0XPR36roSZbNH
u11fkVoFXmsE+K209qbn0FhpD28SSVa8d/E6YIUTzz1Ed+S3g2WpirlOyrIneC0EyO9YkR+2tL6H
ysMlUkt46wL+nPgDfBxM3U6jSwDe5/6sKBthK5E3YoBY1SNAl+odm+lttz74Mty/X+RQHniw2wEr
QfPP3TdvfF7A1o5pa/7ZsuQESpHHFToR+JvLwLmK+tG6Rx3FTuIZyZ6CpVSdFnjtDBVPnVO0u8V2
vL1CZDZ0Q+7Fe4fVthX8eBnOtp6AC/noXope54Z7BPg22YHrkRQNkPPW13jO1WA3lAspo/PeW5Sg
DoCd8u32fzyDHHBAbeTn1jyRvaBTVOxAxN7Yw3GVt58oE8PM4yDOQ/dQSvlwN5K5lN/bYViJLimp
UqKDX8jG+Rxc2vqgnB4I7V6Dsuf8M9ZzOWRhydQh9SQTRUVezgWBDCJc/RWHGy0iCgicq1YazyRf
jNvVV/Dz4ZJwiQCcdmETc6Pu0FTa7nDhr5+eo149jW33vLeKWwX0ZEi5kag2i9cSIH+kxab8tFYm
mbGKu6/mPJZ0qblC1F2LQdQ8eUP5zgNppRpOZtSCTvHoS9maJN7+rjxjvTyIB358iQGVhyc2wn4c
bJJqq0SSvjdG3xVnWhamcczj3QgOq7raj+rgF/LEjrIeDDuZfSCgHDrNdBNRt9KtZ+dFpIJU+92L
hyE70oKJjOi7LY7eUbcF9HSKvi/Xojo+0UGQVESBpsD+EEZb6F84QACqd0Qm0bU38rnvldMxGc7y
RdI2MhMhDjq1FRsTAz/my/H+gKLna9gaLiU4uhYVFJcuHV9PZaa3BnA5kz5q6+38yKBrb0gaIzKb
nWhKlbhM0CEN+lLdIPaUikw3A+fnsc1ZE73UPk2GomkgJTiJduQ4DLWqKNcyLKixlTtQwaAX40Y7
IVfx4cIY80wy0Rlp4un/4OF6nTy8He0PQh2rpDPOKB5hvQVJ4dTrc3VikoZjvN8T3CtVSPm9NO9P
oGGB+ZdJSD4ZlmcvKpLP9wig8AuyXshxzAXFsAp7u5MGZlNNYxwBTSQ2f+x5+59KhGZVkurc+++0
O3Xr4ArFoDmxYDKxJWQqK4N4HeM8bCVvyfNBXg8ZseUNzOJeBjcwksDt7MjS0/33RoSDg7dNW0WO
sdpJZlRKMxA5P/7YW5WRhTwZo6tfsTVIyzZ+J9hOLtp0AxH4X254cWD8jk27S6CZu2i1zH79HSFp
Q7a4OQF8wfqPeB6hoCFhTFsRvdR+z1zhTSIcrPspRkTzgTDn064pEv1nocXQpMiJONNFcwJFitRJ
8l+meuVVcPZuM4IRPrFan5+QiZ+0/lzVA9cvq1OgSOVFsE6C0YpjdykKVy+I1piKHGXTnM8omgEQ
eZMJNHOSG/IFv0XG+qE1BMs+uoP788Q+cexibsT5cBaCEHxvzZUamWzpWB8cljKA7MshnB/9v2I8
Lo2JsDrdvVFdCj5OENCBGhHjF9JngP2Cxp6iRVxxDrc9oX0BoKamMVhTSwv87Wn0xLWQ0MS17twM
4E1cKhqw7Xb33lbySYpUoBDLfDEgxBLCajlEW1J57mrLiX9A/r58wvozzwG9vlqED69A2joYpaQ9
+A702j/X7YzeeaMU/x4f2z85iiRV5AhfbFdMJQwb6mlm+V/wFcGgCO6dU+DKtbl8xe5a50U4XHUK
u9J9NRh5DeWhjYtJCUzjczbRh1avgb9Lxdgl2iVYhkcb7LsAfWfB7axUj2tFRCQfpN/hOtg52eLc
mcUMevtJnlopYNpj1vGtxN0+mZMt9Aot5ojzL3fpfJnm8yQ7R1Wc4uuPRy+XyVj7wqLlwUtbCLDS
g8YWoAjx8PVB3/LFWAWOlOhxHx7oCk+94oRnfvxDthrOznuNH7XUkrX5E3UoUGT7lg9HPSDk0g9z
w33XHN+dFi0UTPc9yxwGPJU0uzPKEE+9Lrj8Fpqrb5Wz5zZ2yr9EFMzMaC+rUpJSTBYLmaqcKlwL
czP8NzugU0EwWxwdrXI6OQT+rJyM3Tyy23GPBaRp8ijdmAtTzuJlGKwnkWK1bFkoyi3IZBMTpRmA
pFSUwxIRrPYExYTswaUo6frPZLF4eIwPvOERUnLx8rCMNTCiH2jxszphof+EyZLBHYAwhxLBEyOZ
q/NpmGvWmCdP7WdN9Bn7+CwYyJb7Iy3D49+IYay5w380DUjpwVF+6521VHIY69iJgyhxTcZo/Pde
YPP8yzwEEjYFq4wYnBNvGVv+zYetiMzdc+y+cnFYZrFd8i4JOvl5hjAxkbPqY0IPDrje2MRWKYY5
+aMr7DP3oXpDbJO4OrkkD3MXjWpLDgbQd52n300l3g+j29kaAovn116Hhg+WFHMMO9BzXg1lqepF
nTeH1UfhSBAcIutzeK1EjiYwvCxDCi49XcIAFmEaCf2SkGF54tWGyCwbNBIkFEGskudNWgxLmDsK
RDM8cNCN9tLQwXaB8SywL7NQ5kvm1y7E4t4AtTunjhsst9XIxArDgdVMgVkJAnqSf22/+S2KI6nj
O64MJMumexeoTKmf0cQwCp2n9BlHJBG4bGKWzTFhpR0yPSaUSWTt3eKzTrjys6FXXcK1AuPNSYq7
VXl++19dDQVl/dsGE99MRa2E2tH9K9l01YF50vSagy/ugZBhhFP6jn6g14yaFRbNexfGrCMxxBMm
lloP657/YDxdaRM3mK/pCsk3XqLuIwQunnmJRreshd1mFmI9iybCnTp0IgVivWMnIQhoiDNZ7GO7
9HWtM7wVQppUoZGUB3KLcaLCPh9Heu+m3ZJSJ4v7LYJgeGhVnEmIouK8wAXnI2jTmVbj6m4/YbAN
Nlutvfydp0q8oeuU1trYi09j9Nc0Kky9EoquDb7lchZ0gKfREjD28e0FCKChOXSlZe4r6feFhYSU
HGTopG1iDWS+J7sfHQMwSHGBHUTU6i3VFKMpYf/pduOZLbb3AJJdHxocypwaiobcSGdiypQt2ag1
h/60uytc+zdPr+NhEk0/HfsIj9U0MF+UmF+w75HoyEjGdzvOjj4G8gvP6Fybb7+N/nVi/Ox5NEvI
lV3TQSdaH+aIOowBkpJFI9oGc1yoG4C5mGqUbZvMoGGC2X1YrgzKXGp/UUey3oFiDZfnhP+IJqcm
iZVx7GlXrPskwvAwg4U6HDiwuty3fseqksbKQ4FyiHvr/2tnG6vUCOWFab0jJxpoI+pwl83G0BUy
wMCwoxICZppuAEZHGi6OYXF80XvwCy+fkw99ArlPqgtFRSbj4XpHL+D3IjvM++TL5bTxK4DZDIwl
NguF2WGpzkD53szSsdx7CxnsML5lajC3DnDf8CcNaYh3wauUIULT8HN2zy5pk4MLQrCrOVqblAsL
C1TyUUx6ojL2ew+YNIGR6YqTL2ymnQD+B/5gxXaK1duxmvDAjaAhHskirRNVAFJNAiNNj2IfxlbP
iFPchrzMMIcneb4yUfxQ2rR3GAejv/WMELNXAzOBKqbPqj+ONDP9Wd+Fy94FVA58JFZWHT7eUT/9
7X+KKD3b2AHQjCMyQBqta8U+iFHP8XcXr86xeI4Xhn67I2AG1P5A0x9tJuK86f8m3ELTjXfHL9k9
w3Q+8T2HxAi+D0J4kSWMUCUExZFiDLnTJOOc7GgMWJkrqd9DXdMYK+GI7tl90XxFW9P9kEXcje78
nvl8X0QuP0MfbntV7V+6bP+yhIzGnjh0kXW4Dl+/BpldRCik8q6/5ZvfAIVoxGyKxAcBj+FXCYZw
GBnsH6Og7Z6DENJVaVDUswqrUbXWrKVyVp6ozARIxa2APQdkDpzgZDuvgOhx4TPEPo2Fzztxmzco
CTeszs/DqFEP+YdxkqA3Lxzfehj8K9iNUJAjqnlpn6IKMzZjgQ9ddFL1haCF9iHMIxvzmYpviw8V
CTr/WvZBuDGMvBlpvtYjY2ncnO1UzMQxyKZPVYCmWxVeNoBC4UhEoqxHH+Jmqc1sjyisAa4MLSp4
+KpQahyKUrYto7C8ndK7rQNOoJsQPv9swzrCJBbWT2kaVApI92M8M6swxZcnBHhqQKxJ6WFCA87T
DhtVEDXOLhDY+pcqamLsF4ytJ1qtiowzfjb/WrlzRDG6DIrqAXMJntttXwhNZoocaE8OEAG53mH0
mnvDKMK2+ipwM3C07l8KG9bec50DOFtuwuc5Xqg0rxmPToe8CGihngYtnipK4rEQx5p0/J9BdPz/
DWG8cIz7a8Cz5HeoY7So8Oa9k1m11E25zUdeYVjZhfsla5XJUyunCmahv/2x2DD9NtZBmLq3IaIq
Su+PdpZBK2nSAf4E7+oLZqJawjnHVk9vKgEiw/Ursw7IMj4qPlLYw/k4k1cjKsd2QP2uczNFkL1x
ffJ9D4nYMRpGwJTcxBJgvszZnQB0B6mTnJs+ytizI39dNfkMiNA2m6ahV7X2xFpvw5DucsyqSN5k
YoTx6k1nn/1LD1esW/qHrwS9D0yUHw8Yy7n/9gB/GTp4ikdDRHNx/xo2PbhGYKb3sO/0nhNA3jWp
5fTZpgujo5gsuVfiHZDJMpqmAiuT3F/F9AiQcJMWoygF6LiZSAAcHM89M2mjEEhdh4a0acKYl/OI
eQVuEMikFJiLIpzfRZwjWD+Kr/kwattPhCBdDbAldjXjEjaqgbc7zbr6a/maB6Q0Z7YUjCFVT4Ym
tbndRuyvjw0toaBji2X1fGJDMH/N4N5PRoHa0wUIQyFUo0JG69O9RXDAx7uKw+3Z85waTpGaIJc6
ep/NjGQElvmOI6rdea+9U5EmKKaLnDJIwCv0hS0l9MsezRkz93urccVj4oEcQHQ6xXap9Bp/wYLr
BuAxnCpqEYJo2VhVEHWGwMsuUtrEmLWcjmnoTAkCN3O+6kiD/GpZt2k7mPp7Khd7jIOHEkmIuSTg
0yzz8ozrZqW+dvGwdnkYxoOjgP1ieflqDZx9D3yGIyWJ8EgJp+nP7jN5Htg7CwdVLH3h5Z0s26dn
128w7wO/LRqdl5vUX9PKFoBeNyv0wRM5AXIJnE/PyYeCOef6xxqEm53qf5SgCezfGwsZcmbwBT0V
0IP0E9wtrczqb0qbOpm2Xo28zIPGlvAO0+IhroMXnrgC0yFnLpCTD8aLdLw1XfSdNBDHe0mSKeBa
8EEIskJgjgkZ08BKKMIQS9kCqrasp++sy9OYwW9sDWdZQw9CTkkcetLzOfEJUu2gEFRI1wMABihR
7eWih5w2xkE/HIVqowqft/xzxqrYPuMxyW8+CwiX9yIKFhNO2+20E0z/bLYV9DbeuPTHQUFx93pr
SuB4as4NUl0cevc1S3KnJVVZit5U4qPAcpoYvuHf5Ng2nviilxYl8LJ+7byihlLZi4iDVLGIwDe6
auM1ozdXs2mie/3R9+4GyHsvitdPr2oNJrfgTAe6GXu4TZ6HU/+9nOyheoVr7TSBcfhRJ9Rz92x0
yOUsvg5J+i52otFv0gVomu/PkhsPyTvU4eedunyfN3PMSwSwV2fmhxzN/v9Q+8WbeTDamy/eH29e
tenkNh2VwbYWzRXe+fog9ZuXn9/PLq4fvtXIdC4PtR0sx4Fthvtz6qJGmQkyGBuGwePbtPBF8UOz
TA9WxECsQhM3CHKglRvLMeWEDLjfbGOFzJKfpJXtOgYLQKXeYUhl5w7XSbBVNXeD3nqevh7m2cRY
S8zAdhZrgcIE1d49BP37qSLK3kBeU5CSXO9Tpn8/rRi8nPdN/0LzVHZuSLJk+MHBXmZj5AyGH+2Q
uiJJRtUuJs/Njl8WEfrNyfDfRmBZxpiTXAxYjOMC1PHrvcppzq7pexy557S64CVUXwIHYdmquXuX
iXJTViRWE2PlhNWMiCv0a3d5lYaNF6YVFRuUmxxrjKXqGjsZ1BWKgaKixCq4U8MI9BNQXUhhVoIW
YtpgjM70s9oW4qNdn3rnd763Mi0kK12s0xRmGVHxNAVkttbWcOUF7zrwmexU2ihXOWJwN6BfYC0c
w4BYIuNwrPQqFSzb+flNtwHOuLrmAiGFlQ4kF5ZL12ty934766wpm7A6Woh/hNIeK0TukcY3FkPg
sH+EelBmwITFY2bv3Aut/TqSO7SwdBU8B1mcPy30vJwkfl/pc49aMLjJ5G4Vnw1ToCCjy+CyeWyz
nwSNweM4Et3TGzrB68Br0BL1y2leEiAFHL7vSGk1owJFCb+QQZkBq350jCEscvye9iGAjHsLOY/5
V8az9aR13vAAgEmk+z9FV4GKyzh39Fqrl8rcd9varTRCy6CMR+lUa5POCQQcKdhBoxkI/gdF+vpY
BrRXfXTU4bi0RdI3WrPY6dp/uZ3eS0nX8bQzKG36XGKAldmuLi1zQVpT7EOYr7Y3hDqvnVAVr3T2
bN0oPHIKZ6Mxghai9/plCCVXAV0tpG3Zs2gVLieMXwapWhpYWPOtoLwva2+MpNFUaM0s8/P+kDSg
gQpCgABs6kBWXvHp7fRXiB81K2nZhtV/mBn2WBp18xTRjS5pvlnMadmu9s+Rcxh7Pj1OBiQvMiQj
+hlxnd80ZEYXjNniMytoXxUM+gylNGBsW4dg40yXZKIWcHxZN4qL6yb1FM3ikC6m562L8L37Ut9X
Z6a3dsJ9uuYAxGdlf1kafPyesqon2nuC8Yvvw7Xjh9Zwks+MgXXs7P6lH7sM0Hp+FEjRVknxkLZY
hnMvjEK8zNrMisL2r3NMkc14aNMRHxW5B1t7MyLzudoqgZMDChICTZBrSrJAF+AN+ZIPysECAx8g
Ewzgyp+KCCpURHEK/5m9UmJSnaoZVxVjDGPcSy1SBAdvjrvn+O0Q3+d15p30mGnxT6IyE9AvT5Nf
8/l6UwM4oFbib2+tVZuRhj3jAvqFjAgMkizH0NMwVGjULFOHpKvCKmQafIpHKCKuintndoEZff5H
tLiJz/n8/Ceoi9XC8hzd/LmSzHZGCMwukNmpf9akiCipyqF5P8TAf6UffNwGBUlU2XLUQkLiQ/Mq
7WOiiem5TJeaOjwFsXO8M9cAfGx+MM1vbdOZgKpPjFoAPgL3elgMHO+zHxlxKzof2I85wN9jPZWc
8hMUwHDlUVjX0xHOl+d57uThVU2o/fbtCaFoI3WUMK9GfrLs8ft3QmxWvbicdmK+HK4O0AHgee3o
PbFaKTW/tZzyhEqTuzXvyW744u4xZ/CbBOM3Jh53azDPiEKUZ0O0Aqu/QPinXaz9W//g/N5hgIkX
yR2K+PDXgogVNg7vlz25ITKGlV7KYoSiKlQVyx4OTctNkhOqiikwf8s6XCt8ixkBzcsjAwgiliD2
K7YbjMSqoKHoo4sRvjq8Zim3sKk328h4M8UIC0kb0ASI0Dgwqtxa0Rm58amCKXWbzc/W/KaQQMpB
H/dCQNscH9m/OmkAWnURYMJVK8GcWIscdAnAz4y+fcpng/YRxI9P+jEB0kiJshpn4Us/6vVrUfk0
LjCJXMlM6rusi5P9763ukt07q4ypUBpjwKgy/YCxJbHDmCRjcmbztjiV+QIlKo3HxoCSYH0hdwo7
R/CEsH9LcJconu3784+Y2OuIOTP/69NDWUnCKaXHBn9+cFHwdoG+mLXTHItNtFxCMlUJtOMZdUdE
PQoZk+j3kTEiD/YPMO6XWo/ALkelQ1kLmFsnhHXOv7fztUWjYZU2hV/SkauD1GCv7helavI955jK
FCR2l9MBDYtmvhE+MrFDEPrOvCE77bbXTrDXPjpqAZnLKym5LSFlEgp4iyHQfM/QQbvWzruvFatZ
K5tn6AODsVw+3UBM6Mqig4yTL2IcH+N82t4zwDXBmK8PmgTV8vuJ4cmNSgeDaVOCRRNYOg+KnLC4
SV1FXU5frWzXx3SOIAHWh/SSld99GfpmpRxMV/vfvlTR71S01aQzmakLntH2OV9gEV9z+NuV5YgD
+f7ukk7MCQWKP4Tv48ugX4E532opigkpjpLqOPhkEmTFgOpfj31iECpEecuxRcrnU6DfopiFCMcy
EGBbUffjiWBg0nwvMq0+PsZdSByYzq3N4lPy5lflFBAV6rMnJnGEr3Wo6DVNcosAXcn4nXlBA5ZN
kYMkqpMU/gM624mSHeX1xw2U+Kp3EQg7+3PX30K0dMDaaHrVL3YU8RvVineBUOrwDZQME6RWM+s2
j/VIiliSuUpw37NMUl3dmTukv6yrUgzxcMQg2byZtDBTtenaDy90LEvXBjX7NaHKrjYnltKCSkWc
JKdGmik8t0og8C1kDZfN2WaMm/Gz+T+7btFXJpzhxtVKN4LYTdk/2oxE1fhlc8d2RIkp+zSAJC+6
p6qqRHlyLFdjvfr4ETifRKxKxrttBXD7JNbL3/LWApB8G+KCC86/CgBmW3A1ci/3/jSeOzzt2/z0
F4/8TfTKP5tS9vSrk1IMtnUhKrxgFrlZv9imRjmlIYgmbQzClaEYRojXa8x8wNy7cadPhawTBssG
XKVDLAk8WC8mLU8hgZLUm5oyqBjdBu6nZ7VOwzM02bfis/+0IYuc0xarW5etXjmwgFE9WjID4lLj
7F6yU09ms3DuH79Yk9VSKyq1zsu4svoZVSRHBrwCua673/W0kcyXwnwHY0OPZVkoYre6qYoUTpdL
wx+BO4ys8grHykTzwnPsF4CQXmB5Xoya47tk7gbXQfmRdiSO/XvyuKOJvlfmKvio/UnpdNbta0J1
hBGytGB61rbViHoARi6qLulQ4BHcMo0ALAwrAMgXG0OYL04pwzpuqO+BDSWASrFdvA49JRGxtsG3
gs8znNTpcHfriYef84Et7oVRqh7/gea4OBUWE9D182bFfoURc+Ib/d5EFpdwLMl4tSy0QF6g5XGH
mRLlVJo/VB91Xl2LEG3ry7Tx4MIhlTnS5VE/hALce9c9ODU8q3VqrjPtU5JkC6nKnItSdfsWmooh
zzY1YNDBxQa5qAO2g/fNKuOILBCeYGQ2iCG7+rXoQoF1ra9kDbD3cwDkS/0Gowf3QQNen6Wk/WbI
t1K1nh89ZK6Z2EfhA3G19urvWi1fitpp2s3qTiEvDHzPfmN9BtjDc3Rh0AN1eAhMXiE7hVl4hCBc
qi7Jn5XM6MD91jCxux/50VZ82qAVBe/4QB6FzDJB3VAuh1ussZfalYxTYz6GRZiyGqgb4H/oj6h6
VDNx/y/6yaiLwAEHi4ndJ2vysPYXzGB4l6WqSOflvTXecymKnL4/blaL1fqFiD7GgE/acXYlcP6T
Q5oRJaZWcca795iBuDtJyi5rYLNNlKZH9XeF/Q3J0XfaNzldlVyBC3maioS94ZCaMG3ntGlZHcTs
XuhydiESF106hV3tmYZoke2WjsPqigibrAq5yhms7LPcD/Jo689iBkXUs8230TAfZI8MZy7pyY39
KfcnhSjHtVA8oUOlYYMZf3/QH/48q65/9nCjTa1Jsp4DhQ0cRoLpnWf/hWzKKdrR7bv2tsWQZMh5
qiPPU0LJodhtAs1PF7bzdX3bzxcXhQqfjMgdpxjriOAcp4d+SaKwclJaLEudGsEWHylTxQ0+ehxc
1eZlDuVjcJem5NxcqcdJmtjla3f/lpM7hvs4xuAKIX+kgQLjpzrK8WFPGLg3t/YDtKidYE2YTACl
vrvjyyyewhANi7I8PffdubzcUgR2SKy2ySinCyqMCmpFnrpzAyEcJA46AGj6h+vt4xPNZBDs7vfD
KWstbF30vEiDN30/kvDaKqmU9o7LHrgcmsSkxngMVP8hzC+zUyGaxx16NCgfPtpVi41owLdS+JF0
Fw2buQwCldmbQiBMVKkgwi+l64D56Dg2GRX0GhRBYGGIC3NnlcLXEPzpMKSHzBXTrpvcqaYVLyFc
RpkR5lWbob2TWNgmwYj/UeerGctGaprH71muRajLf7y6X9l4vxU3t6ppKjd87AoX5F93GNc4Bher
wRk7LgcMGVIN1AWDO/hlfEBsP6mgWzINeFZjRWF6qjELJf4zFJRM2nWpZUtoeo7zLXx3Aso9GRHz
5yT9c4oU7dYp4/on1kgXXBsZR+Au+ZpIQ0/BiTUovnRKHSUxZTfAUfyDSeGt/Xkh1sU5sfInGXJj
0zRfgY+ww8kcyvU3+1Rf8f2+kEE0IthR0OUuygHVN7h30dtJ+SJzl16RmAAAquzTlVkPf1ZRuCSF
sDiw+z0TvhoVmzIDBCrNS/fJbxbWVQyXmpPb5GLuGSjeGA8M/KVa4m6NXrkmW6rGoz3uLrdcWv6W
B5n+rRt85AKIrUf5vJY9KdPyDFPHFYzAjBWwWSrp9DZe804DKoYYZyr6gHgWLdxdyNJTFBxJb9Kw
Um30SpF3cuebr4Gi8f5V/uYs2c2faZElRq0prxJRia1dHavkG6wX9QRHgSZZHRTFKUnkEomJRZzc
DRqNy5ZoGLFAyEMqmqXCG5Om+sfU6wf8ZjvekRtfJLtsMCfAWqDWoLFkpptl7fwqYkYCdBxaXVRi
s3WGJwA91q/HZbxFsSxg+ZK/2c0rP0AlI8SjpRDLtX/Coxz3RQ3pG4U08aUQmB5S4dfQmpB3Vycz
sP5KoqGMVeXcMMpKJQBltbrBKecTl9SJboEdDR80UnQD9hIDwd4Ji/SJfr+DO9nv4KVAk6OOq9tw
fZh30x8zoCB964iV/7AA+q8AD9MPCpRpadJruL2bBghQaM20aY/FOEAVhAGU+U3o4MtzXq4wobMS
yp+o6gaWOcswLBHiaPlumyPJduKREtejYwYEnBDPnskw5llHx/Xs37GocyOGFSJHQQcV8eGB1TWo
PWzL6/Cqrkp5sgIjppT1H3kqZB4f4ipcxOGPQnMQ0QvbgawhPIziC4AuqCA8zZRZ47BVrvDWRZ+k
H+D8BJXeypDVdw+HXFZVZMAm+ty2o7UkfXARDQUpBAjygmVyzEFBZEsV3dT0PLxv0eBpd9tU8NHI
Rnj87lqGtZvkHEqfvVkMEcKT5V0Xnj9eLRRE59Tnjt0Lykv3xKZxJhJs0W81Fl2s6bSLzhWTFrQ5
dCUZcHINcMziKlZCjHIvMgeZ+IHcC2uMXxqOL4ojZ5wdVLqWwvyiLOQly4TS/GK8L/iqIu7s93TA
V96MbTXJIvIVhmrDiKyO1i7cb7yfHMqALoMd1HlAg9PUdZ5Zj1qINGnLMPVaDBa5AEkGwEg66FZn
QANYpMwgVl3H/FvwSKMvF0nsvr23+17ZTQ6XjLFOsBj/kQdyaNTjMsO4fByAY2RoYTC3e2vOokSd
b8ug4WiaQ3KmmGtOmGxHt9WH2IpHs75x25j72NxW3EHmqCnS4AIf+4ydki0NNUncDSbeBFuYifl1
KRJTlU/5xfLBsIIQBSSCBis3Vg7mDfJjTfD5HJj8dVW01mVrA2gT7Yr1viabkrWRbUAcOI99Vboi
ZBj0L6warF500epjFEOEFE48goEzBUg7R2wZhJGYhy5OS13ohLUHKXXsq6R6jBNlrcPmr1Fy8AbT
0PIQPll0I10PaWq6y2KO+HjxNi6PhoHRJYaO9FdC7BHnB0/9At8jY+Z5fPWU8c1Q6HTYlgAmlCIp
hOhk1qMr6+aFyFfnJRDhH0vzIxHJOZ1qs/urkAKn8yIb7FavBjWJyok/FHktCMoYjfYO20X3RT1M
w++yvDYg0M5c5y2itFDgwd4SxteF78w4qtxFAeMlWccJfceRJGGA6DI2SZtMIZqaq/gk/HR66ey0
iUQCGa993SI7YpnEd7Fgr0sF8dOwVhy68VmV1yfQgz3sErYF4T7T4ccRAnxaC7KwJ5zBcYF9QKYM
yzHVuv43cubq7UAYdvoIPtIMAxlkZsB1QFuDKPh1eGPppsl7PQ/4QdENGifk+SQSiF/uRlEyI1Ik
uLewfHFdPucu0WL+Q4WUxekjcoviUFA11XHWeGr22xwjkw1x7WK7A8YYgwtNTpLO1A+cDLL3GvZC
B9Y0288m2wgbydXz9xwiKFd14hu1XncVC3iFf9lJm4HMfOr5H8OPSqaMaj/+VUhp0tIQ6AAjebCi
EvemZtEz4w8/Nf8Nbv4jU+v8uaguV9CMGTF70J6HVkA+g7SUEW7gx41ikfbnSpW9Z5EL8uMtJWVA
0fB2O+Tfy2crGCMnnQGbI8QcPAypUSTTBi7UhG5ulBMq5Yn3k16rwOq5m1TP006VsEAMRY8lSMpf
0XG1XYKbBCC2ZAxiwaSFl4vcUVRnn0AFXMrZUMnmTRAiws0fkjgt/HAi1AelPxXbAC9Gbyba2UlO
+N5uvIBWalPfAxIjZuv5Jc9EeCPhxjhKAhov/i65iPXUKrxpc/YSCekN3kUHr+yAWyy83lvV/aNH
t3H9iF+1DwZBSZ7NkbO27wDFFa8VbZDKfmNHReru7UbTZgbWFIZZfXlGuDqRYz6XWmR8FyTZnq6f
TVCnniBMiYdYzRSXFpJCV+yjGLpRYifJUy8IgWtcDBgmUk9H8cdc8usz69a0+rFUOuEXUewuhJoZ
THCRA0+6nEcJjstr1GC7rmnWJ77DEfhdDY6Cs7/0c2IqrkFtwgwQ2dQaEvkb9BlfIwc7FUpk0v0N
HZycho8mQEIviF3rQwn8OuJPluq0ZhTkGpcD6NB4uVQnXbn4jtHKtyMm4WsGirXFUaTXb6blXRM9
s96TDL6tm54fIbOcvKcyLkXgtyx2CNbQ3Dsy/n8RmckpnHwjsz0OuUPuHazsBoF3dws2nMdcyDQ0
NZKoWiX1f+dFQfhtl1V5jJ2Uqt0HEodIUNXlYjNJ/zvAyvptRYD/38zVKqm5N9dgS7OKT8zfDEAI
4lFKoKBWRfJ5OnjqqNY/KlHq+JMy3leNPjynSCifLuZ4ojqSPiTe3pwxMddwqiJCCJYHt2E8LmoP
85Cyxix7CaE0HPbIdGYG4T4yrLR68amUaYfr4n50XR5gMIiiW19MpcCICY5VGUyhFXuIsn8lQZl9
8QJfMDKVLCYEnSnRO10Xsx7K0tZ9qPrhwLfscv+yR8ptPTSefBpBLQHwhSSC0DJt3raWWI0PbE2C
gWmJziqcVcGDnRMUkHaEd1/oL/z0L1LUW9liJKpAvvW5kHQ6CEafmu9upmh28o2abkMZpCvJG87j
U8pqQGj/ji3a3pAlIQAkAkY7gxw01y9jg5hgDKzxxdxhUUzFgOJODpUiS42pz+e0vkMnS9nM9Ov/
37JfXZjXZJUvHO24vi7z0XtXJUbxXYS6DJtzFnHlCzl9hPOYwMhfrLOS1/fEHbXOBkMRYXPDx+2J
zm16UNy2Lt6lFEl+p3xlWWob9Tt1A/5SE4n/wY5keTm7NAHjCExq2orG72o7Zgh2pbuImWQa9aP8
emOBMUiyg+M7C2+PN+Von0E6WGJAnf0HKdJHoVLoCUToUM3fBfOWAmdGbuQJVLYiQ7mDDOdPMrWh
97yq4yuj/nQpdDTCxGTNs1Bo77OMhKR8fXUnGDOyet1I1tlBPPVdzlS2KHbbG+fTR2Vn2zeYq+q0
4iVu1lSo22DF/tkEflONIA73OYltCscK7xlhYqtF4bAhHr9RQy5mqJl9WaUBqU5Lvs2AvAhWipgO
94/KnmpfEDJDnb4J6xTgPvF+hOMbzu1qUT6gLkd5sKXoREfiZcHQfaHeyL4NqTUXgDzlcg62I7jV
LU5hCj7paCXJwdDulILNx+Pw19X64cpgleDbDbiAdf4pe0UxsJERn0qeykdLCuaz+UUUFtC6AZdw
cEjZrJVODzQcsUwlokCZ372GBPQJtb6+VIyqxaUJO3FvuDhvj8cQL5C7YEWscwcLDuF4I36xuzjk
OmTsuyfxoaaH97yGd4y6DOUi9hECMRwdNW3Crn5D8KkrAEFILVmA83A+fX5lfdvJvBRdD17Iz2aI
l0TGrkrbh9NkrY6C0PnUWJ2EYLLYK9TNuWNyGTBXaa5PuxpOwuuSRqAkI8zjD8I0ZLM6G1enRTLC
BGNTZZn82RT1u7cwcuBuDCs3nfU7CWHQTbExMQOtxmOnsfKSU13R5jLz2hVv8XUJURzopLJfVPQi
EDQ9bebQ5VKQzuI5ELWiDT0UERM+7CWeRcQE4kwRHVOO96mryQhS/rtJlDfLPNUlIu2ZN/fb2OEx
oDUAaeuCUa1KhhLr8yBM3TDs0WjWY10JWtmu/UzV0niM8se/4srcI/qgCeISlMWNtQz0DNgjBLpa
ygj7fbADhA+sk6i6BC/fPrlYo/rtJYFwDV9+loLJp28+tBZZmw9s/6QXaGMfxKVBAo8dHGg3t67w
xzIL/hzzbdjYfSx4C0UIFEUGmYj6fUS9+IWfZFPtrzQgvYSgdOlkOzZoP9b+cY9feAqOJPg7B7MD
UuztWvxT3edT4z4tH/dCi5z4O0eqnNJ64v5bCSLyL2k1vkEfhCgj6br4A8wZIHPxy2HFdncGa3IN
vQjRuWBj5qwihSTpVHX5SiVTiwb0ymIXdnt031bkkB75Ax2HeR/kZMk/aMF2aFobshnIfvFhlxpI
Daa15kriKrkvwwTZiCqC1ynd5FRRt+u76/WiIi82rcKU8+if34rtlKJlJ3aDJPahW3FUR4XVonBA
IMHvcHBjAHc9uQboRz3VlU0IuXr7N8kgdVL8U6g886NLCb2bzYChQ1PEquFkvBA2bEcBS0wgwycf
IiQYGwu79a31nK2D72Nluo4O/UKO+k9Kz5EAQubpoCmjEJBeTY2tE/HYM/B92RVXcWGUhL0378G8
wBZ61SZca3PWsY/U8KYcBiQ3R6iymDGX5m2K/t+1Op3mX1JROGpQn1crosgeyEnUCEgRddQ/zuJX
I+B1PTR6ggNIamYsgwMux5tAqRcS3Xg0HMXcWRn0k6uN4bZC5iZG5sC6w38hpckHAkiGAS5JcC5z
7kkjSMvHpz9Av4tqFe/HbXc9Tfy7L2yB6PflBtZAJvyoWub7RoxoOr/uZ8U4crpy3YI4A3CXrjlv
xFv6NUeevrHEO7DY2rxZuCXZTIuMsS6iYdcdAhIo9LO1uki3hFxjVD6dUMb+viPDbYoinhFcdqXp
XkSFMwHmO9OsnDkbqXF9kvNlIfWaO/iJfJvsEC52rcz1Y18o1vmzdoIA9In6e4g1Y10GZYkwc4tS
MsykthC+sPCqmPFlopgSiI+rEnYBjsW6XpVF+7aM1l3SvXutCPErTPsdYK5UAEDPMNORW+7q1tZA
TFP3w6RdA+2pLo7X6ulJorgV2QlOEgcsj5f8D7ebVdBPa16vcXMhmHo4Mn110F0Xc1I3lEmqLnbo
ncpkH/Ypt7kxX6cwmjOyYfs2OFxOeWxrXgRjZ78GptlScNG7JrmYfRSD9rJuppdOklnlF92CF+ex
W0L4Pt4dd0wsMK4ZlLcmnskmowuHH0Th/NESCASYzlaoPit5MqUvJp3y2Az5B42lt7P0QsGyDMNA
kLfyGgpAmaZ0WCJYyww1oDtY4vbP408tTnVL8+YmrfiMR3Bqf+6J1sZsTfR1PGfEqhqWHtBaGRMs
JzveTkSADX8ARXB3YsBwR/M5FgEY8onos/Aq9ET4dD6sm5WKCgpX98+ixnFbQAx7cG6G19LoP9OL
0fce4HKLYqXLj80AATXB0Su1C922jM/9f/m7SOBNhjT2pCILscb5d44+yiPA1iB1g6ptDwVY0oIu
Okf0RCBP2bfJUh9C5PEWKU7gMIQdN8h83ZyrYxrCPSvpZyiv12Gd8LlX1VSwbJ4gCwD/G71xUD/U
exKr45AR2p3ZJ/UyjHOkh/CZtUEpE/UtGgAeBSfYBV4cfSoXMsHVAsXAOunCcx3dVl0FEMvQQOPU
/FYrpiLJF4h6WxowVqlVLXgZ86h5aJOCk+2ZN+wqZJ65vd/n0cCk0rIYJo0W+PKOlV2lgMwzrLN2
xsTuycL5+hgBoePBFizUuGrBQOonhymu6klXE3eHoc6O2FNuA2e34AzhJM//s7n4DuuMeIo2T4vE
5ve2a0vnzZ3HTeXcatoc0iSdYSB1O+Zx3Rln3xbA98oWdIpCoOpOqdX0zozWdj7mHM0vgXR4vF4g
LeQaaFUydJtTzfsFGe3I1ImPOL459aziegfLLIHOsMBfJEC9cu/DXsSbZvPGGPFRvxSJdu4k7pRc
oMgOs9nhMGuUTR9j/VkW9RCLcZDeSMP+wgjXPPbyN0WAmCqFjlnrUciQobHxeQqQ+UJqhrg6gfpr
9Lf1RbheiqhX7HHbyqESE4Dppkoccxhf9uV1ukILhI0jCXAuIQKqxivvAcmUTC/t8pPoYzMPxhLl
uEqJM36HGLG1f9U3YWeNx23Lsd6GnopX/YMRNLiOaTy3V5VbWYWRg9gdcuHGCfgZlnK7xBCns3RJ
42XUGzOGTioNeE477D5GKTdx0ObM91BT8k7ahb2hgG6nFYvTLpI/fj1lhFxjx19iNBQGs8xoOInS
Sj51uq3d8WUXEjPZaBsLrP0dEDBWx498EQEvtWn+feTOJA6BJK9cLH6CnzIth1VUOFYy2e3B9uAv
W9BD5J+vg06yutUwixC1aAg2DX16aJk42MpiigKBl7/eAwa5zdMWMZYjRBPC99lcnGV4Tmm7SHsd
TkdytB8NwGxAOEEnrBxO2Xy6VnvMLdj8YPMRCPThP/AkAbQH+mJ9JGfLe4mmA7mHcwgQti7X8qak
eUbyhEh/EEEi/86QqO5R6haOhKIQL2HZdpS62ZHt7Ts0tUaCFGSVXkZAB41v8ya12TDhr8LK489e
IIyyOa1WD0wSmoqWz+d0FTdMeS5ee9EFd7/tzpw3qiDc50lOtPy5zVNWFaP4zmWLSL9rPQZPVdeh
rX77HWFHMAatTYZYUvtSozzhF9Y9z4OjGFXYHbeySYrAPw4ulg3bWPCHxOPJebaC3uyRjH9Lxa0n
UYSpKrDf9SW72udU5FpBUlzoA/f/fGyGBn9920buuENMysr4ZQwATuQIEjbu9kODUcxvW7E0uw1L
A73n6HJCeDFSfjeFE9tTbQnaByN05X3Bk9KUnOwpFUPM4F12iQ/6guOlVYa1cgA04Knm29JiAhC1
mY8wVwRHiIfukVV4Jf36bbW7udz9xoQsSG8VYUBwzbdRS4flH6OMr0yJ1O4XbdUI88WF2ZSi0pbp
llerPrg8lPagxlhrJmfkyRE9o09VO77jug3uqc5JcwGLorEiTm/RBJLV5ZFKGnio8nUg89v6xuiq
9xSWUrI6QGf04Cvz4pFbvbSSrcBStv41XI1joSJR2lkodQBOqXjL/NtWBumVFenJV/2oArFGxRqG
zCfnuraFQVMSQ54r+137PkI2CocKg/Nh0acbxo2KUo8UJPnKGhTvtzuWQdzTPsZIHmfXPY98k3D2
celd3IM9Rz8VlrcqS7NltYxdWLXz1UegVti/VcEWQgfu7Rr26mHxVlew6CvZCoEY3lUNLmiAdD9O
s5NUwuCWfEvxm/GSfbc4qJcmDlgcal5DTIgYtxY7GVrsO0l6D2AtXe6vtZL9xqFO19nGHu3c38Vk
AfUOZmjNGJ0MqMg/RREga11weVZJac6S8hiL1nbdpxsP0HIyx2+PRDWyBLM9Ulikk6NNuZdqw2Cj
NybYnx2Dds4SjdUG6AUj3VR7X9tk2q6ENXDk4x6lzQLll6hU357vk7+CJhI7l2jTDLKqOs20EcMB
RpM5ccgt7MEMEZ2SV9H0F5AuaxDfZBtz6nKZ00AESRM1wyDAksyjCIKRsKGx5C1AsFQCBT3E++52
q8P+qQI/Ll/KhXW2GG2bFJ8Qkfody930NWjPoX8m4+7XxvIyCS3J0NGhZlNC2+mAKAuYQO2hovoL
yxyFM0MkVmXycgOJSwaRZkd8IvATlip2l491Sn0woRdXl5ZDRT8VE9qoa5hUsYLBoWhfCcKa8gii
2IaHTlrvgD/y1K+MYIeLCZhGZV/UsaLNdf0cVlu7tyNApGsQKZUJytV5ij9HXjJgpj92NPbytrLA
1vy12zs2bseIQoieVgd/GawPZmCbp9N4zT4Ed4OpG3Typ0nNZssARBi2fHWtEHy9Cs/mtsrDwmmr
MDA37GvLj0mu2led+d68bFhYNQRPjGnjZGHKrYmYIaiW4+A8AyQQ+J7IgWPSaAO+nxLPiGMZT9Xi
c0OTt99A3qWPQjl4h5FUoYjebwfod+YLw+1po6wb8BfJW60y1xEUwk2WQpELKO0Q85CQHGALpkPX
gpDkj6ZXlzRSuyQrVTDF1xr41X839IcRy5uD1w8yKPRj9xLxvr/yqn/k5VRt2WLPv9FeBxzLSmAw
SwS+UcKq18ofbpc8RfbPEWD/07/N2ztChfC6K+paBu0s1bTJc4CMbxsOoxIqZKqiplA083QacgCk
xQ71sJVrD/l3laHNmdy/k5AOptYwgSNtTFdNbD8Wqu0JbG8+NS56OKIxSnselb+xy+w0826Td5ke
PtOWJ7in5TF3jwmOwxFibU5MkpTpJKuS78xI0Iln2vkDY+qfq+ym7o4dwNGCVEZJxm8m7a29BIo2
uhbQfnatSYUVsLh0ejajh8yTTVusHkv5s/1FHfk7tRK6McFMBoFMw9DRlQHz7WPE5wsMghu4ttkQ
BDnt98qTi8yVjdOxhgylOSIgZSPN+43ubMRcT355LXkmTXbVEoSnU7rAd3btMaT39/+Vm0UBmztq
CAvbFBjq1S2/yQ1omvZgc7ZPgMvu+KBkc6KENJsCn+bxtJp1Dn4/1/HEqYRtRFWur3hIfqw/r2LL
FW1Y6AqBX5np3GOVCbiE4KQF6x0ylsRDM720kNA7YdIWQ2Xzx7VNgVqsuQlurnLkvMkE91NMBvBX
jrNj6OXYs9p3PMeUkh+uNvG5R0zlmHvE6lBnQYBpic/MhrCfZReH6Vqh0gKLdQEmEd3MfMIFVxx/
IxQnIIEGtj4NqLS74ygrsS85z2FcWpmX1mweFuO1Y1bN/DK1MC7hG6xsLHUsOIJntg0EGQIPHX7R
XWddlUfNtM37OtWOpQIAE9hlORIiZXCFD5fD3jwpBkJmC/W5UToSg+veOrVv1lR3cAs1JR6UEhqj
AYupIFAOek3ihoSFR9GEIrKftd2G0a6TVXIj2eomsNhwWCpp78yqoAs3PALfKuvNinSzxTrXAW6v
e+ALlj8guusMBNu+ijiELy/d6t/gLU6l6meBymQ8qZhM7zfagvs0f3P592V3hqCWVvQVO6J2SCeq
S9nS27FopVLee+lunVIJuemvm9qObyuecGoImrfJZwSpv7oi/wJSDEhREIHMFYLFZZC9sQx1mfKJ
1SuK7HR3emZR7d/Mk255nZp0/k0LgzLM9IfJF90y+ICaSd1lNjbGGa8jbGfbu3o7GTZ4BupjOuDx
Oy04PXkP+3Jfe6YZpZ9kIzSIFBO6xkJ9PXaFNWBm9Pq2YGODhQ+hpalja82qkwJTza9dw4ZTaTU5
OYUcLGgZGjh7jvPHuxeGcv3rEUUAnOv2m2Vj6WcH6g7guOBMveVBrdMSdNOcpdaXM5SFr2zkTnRy
HN8sEiYl7OqkUv79jCaJ13wDZyUipqGiGivZ95AjhOxI0QkT0kFG3mQzVKq0ZIFCDqG3aKtNK0TS
ljcq0R6eyXjZMNzJPpscw51cEZJgMKnP9tayhvYLKQA0iwFSX4UxGj9L7LngltcqHf5ehwq/AuLC
ZHwYTJqlpy0lW9h4xKk6VMCHD1W/COi8NWGP3NL9UizoNTwpyyUrcTVTpcQSa4xqSQUMymy7VbRU
flRnjM0WFmuZ7Y6bJlieTMo8bdj3joJPZiEgMGDhh/UJTbHMxXIPijy1Pdp2rjAYwSRxqIoeYhX/
HU8zfLozAgHNLf/xraWQkVwW1Lvts3Cos8dwIXi8lE4KXiUNQz63r8k8/BoUloa7t83hf3WRC8aN
cMipYzeKejvzq3yzH2+pyIDex/YpKT+/em1iJVkEcT8LlIqbdx9H9fn7uAgTUOVJORjPT6kc92zT
QkjnByYDI7fk4W42O33HzfBd6IH501a5VzuNpvArE5DKPywAYlzK4o5OkPdIHUufZ0FEKH/8gEF5
2+JCLXWUtR7AL3WOB/vkSw2l8CelrsrHWoelWlHgGjsrQC+/pSlhhpRXyQM7TABHOcpb38hmBRJ5
9tDpIbdDmQ2WU3eJ/eZRNCEKSv+eMtGR7EE0NAyb1tB+2FBVnmP8b6qdJabmL6ZTijMWZn+vK/lF
9fLm0Z0tD2vzSE8174OkjG84LwSkyMqHQ0F+ECcilOObRyisWL+laToLP/DeDr0GHy5P1D3OlMk4
99VZQQ0JrQySdPOMl/osgYLLyyndgwe3pRiIKhVc9qBjG+h6s2iNhIjldstKzIOwtVqvrslxYY8c
1JtSZGDrmdQOfAEbhBrIK2aYXHaG0qN80Zqmj7lwM0wVTrdMxDTjdoNr7hzoimTYSghC+M66jCpi
MeKS7iEkU3vi/h3kGvf0eaBSqc2OAM2yPu2IFTJ9uQSWPkLLmVilylQ6Uco9083UJRGHGOL+YYwR
qrJdJjNSIvyDr5YALOlzd3RLWB/yJig+uJAXjxB+oQAYom8ilOHd9V9SiaW+UiR95IWW5Uk43dct
3XjgeahtYjZku0w8mJticyk/1Zxg6t5LQz61IRWGjuRcVXTb1Tp2HuJD5Ggov/j1ugOCUgOg0AeS
G73sAVVsDhn33wRgeGNMQlD71Nn05FDdXmNYa9pnQ4pnTrPPO16eJv7b1ggvD0owCCFuKa2JCG0M
IGHkTZ8kLjgDk7w8nsOLO8OyK+1Uyw+5wwZJIAaq3n9Y7fFc8N3JB2EAoApcyFVP3uXwFh8GfiQI
MoNR1PNJ/XE5TNo07ZZZwgPTM/nGWTbgeflXkefHbAOaUkTawv2YRgY0frTvaIszA/3QaOiu9JCB
8QjSgQXbqnIt2syCPWn298zEEfevLJ0J17hioIf3d0/ETzjcUV4hvforA83lRfZt2r0zitrjkhnp
ISLzDa1YW2gHOUj0KB55M/sffuuEu0/ECOTKhzS13+ruLngh5pw1HBRUiEY5N9T/jlQ4iWq4HT2i
85AaHdrpxdLt2+mzgFq4Iv4Iyx+1JxhDPWm4t/ElubXCAe99IeVY+UjeDh1xtLzNx90OtQT4vewn
aIpNjVMzSPUgME9HwHhIzJhr0/+ON0v+lkR8U491L7xx/Alc8wWPbU3JNpXZg5z1BoiUwxkVSqun
c/bTYhjUf4eipFoYXtg8pUUs5S/tRRH6GXFDFJWmloz0pCNEt1V/B9Hrw7KmIGLN6/hBP6QPKI5u
lZOcj4YU+jLbR/Q9Rh4X3V5VUU+rliumb0tk5hI6RvZxWKYt5bFKZWcCEwfVKog0npnnw1VwrHry
rMt/TloU5vHALdpMojMWyf09knnyJQ/HqMRAgO6hsq43vwTviPk0wfHkfubXreU+7/ghrYqFgnXB
ikolf6WUE/zjz9rr+/Q+A1VfJxI04rHYEsfpHxaKLTOZTzzoZQmIqaaTvl4e9MqehY9A4A9lTCTL
cS/AaklkRIHPQ07T/W53x0KlsKGaorTPDCw5/prXxnxgAB3U1Vr/kgysI6eccLdSYYU31LgOdgXd
jfou+KWUp9DQIH6Jka28DZ/8eKwlcRrzZ2UOMI3eXtQTZpBGPu97iiAQe8Zy2aRn/T+0l4Asc3+4
N4n0NP+QV2nfe9d9HxeHJ5lAsDRIgGzuf8IPougsozNmpX7wjwuuNdOvfOx7b8a6y+raQkI330mw
5L1dPI6O/qDdT07SV1Fi3IiBmiHew+umMlLQdtyhgJ7Xol1Oo7Gp/sDLVxnnRF9gyAhrUChetmiC
bG9EdDMigx0ARp0PXGbVLlRYpn2wzh0XpYbNEJAsJH+F0VrEKgm4NBD/htG2LfowRZGgRaR2NVlM
5CmvCdqVYCznsC5lGqRO6BrO00xXedDy3kiO4xd8wQD6uN22mD+Czwk9smU/BLlD2dk2E3H82VIm
uUItWhhw9WjZImO4tVyEaiWQoLCaEZ+mxbC6ZVNE5D7QTS9UI5fsQ8ctZY4jemGd0AO4PDgup6qY
OIUf2psTErFU+BkT/kfqKCkz9G4fp8QtibCiG9FJIKqEncLXYDtq19smvAPOlvyEXFlOMERRqLYn
Il32M5pVchROzqH1DYAB81nnEGksptSZ80NlEuG81qo/fbCbPPz16A36A+csBB6wFe/PJRLGjhDM
9ZwpFk3Vtn5ghbIaP8BCnBye735/xWCK8CsAITwPpWQuDli9gfupAGgbSVQOcDTygYR77A0X4jDG
1AUJ9eYawuIi4JXuLMmu5m+ZvdabJ6qzi20G+7S9HCH7IzYP5qF65KH4FWnOpeIlHN2iiMD8JPLs
gz972VvhTBvl8bbKdM1742RHn5MvZwEtl9vhk9OMMNufizV13MIEj6yUVmpQKgklAa5zRFB+egpK
gO0i7Mju0KlihMpgPFBUk4wIZv+YSBGQ/XFMPhXRcyK1sxHv3bNySNDhWgcD2IkN4MgkNEmnDx9P
Tb4aWBRjExWA/qUL4ifeDjhBhv2veStm9/X4EKOcm0y/P7BjM1xE7knnvD/iWRZLPoRzDOdXqbxE
9k2gywtT43mKdRxtRAB13KJHMGpjaEdw8IqmJEesMweELjoDm+u9JJWeNYwE1g1Qhw6F0SuXl8SC
fYPfXcxWPnm3/oRIIRItw7n0bxB1iqmtzcOkitLamEWxFjLgrkUUNN+HAX/DCJLiBuv2NABQmx1i
szT2xIzsnlYT0MtRNao0nlGSQfJ6RPVk+lyWgp+vqmW/1HuwqFHx+Y5EU8q43Rs+EzOaDw+vWAED
DbScEBUxpU4lyWCQ2CMGKInwV7Dd2iCCJkMY34lNLwFFxlB3mSiOEA0CZQ8ycO3ed9w/H/qRxp/2
IGf6g5KVPEWVQdOEpT9/xGh82kstsy2qbXATi/T/ELcuroYjbZ58z6Kh53C6ZXEZtRLsdCCCuzOg
i+mqS7FDhH++mObxgb2F0ZtoIVvDBxAwxGifosA7xXCawSa683Cqd8nU+LBILHBP/GnQXA4ulZL6
nD25z/NNzU8MwkPRBASv7tuD1oHMUaTzgPkU54ePhoW2OSfhZQu+K/ue3wlEY/5/AycFxiG+OkUP
b6PfQg66kb6G3MF03cliV+Sjl+RcJiXg+G7BM1XVubPNK7oWAuak02Tivnw7LtqtbuejeD8csAP7
p4WvIwYaSluhcPbSwWhbonf+n8mxb26Ul7qRBjrhbJdtB/nOVMeDpQXvr/jLyVjVlM1OnhTvPLJl
EDXlbW/0koyTz7G2iajpP5Y2s7UTzzdYUJlW+TXLnOsjstN09hpd6lN4T0sKGahq9bx/tKPKkljd
fFNpfoIhGPUPeuXBiwPJvPZDNJ/BKXb2ZE/fOry1Te1yUVE9cSj4/wsXQ28bbp0VABolkvF2E6fv
LGcFPiqTlCJUG542cLlsYKadPueaxl0GouJsPjT/HttuI6j/EzQ1dJrMMvOwcLHHFTxV7QY2aX/z
VfxXCZaniiOx1YydOpGcZGGe07ZbaoJGegI8/uldWIUu3IS+o5aaIuyhEf2gd1TefI8rFAuiXeY1
bBIbviz5XHZu8svoeKdYuheKcKT/Gmebjs87sUd8MuwrlsGjWYUWbyLz2dAJKPRvbs038I9J1g4J
ap1NmYzwNgusJfhrPdwcqvlCucHNIZge83dfyXezFXayJcAjGapHNxHoiY+gbSnQjWCH5t+CwhDu
Hq0vkH5W7rl5zJkuA0SHtJQRp4IQBcmXF2dKlIDJCuADw2C6dAp/YQoffAbkembxZbdmJ8gW9bYN
t+zDkB5XjCXW9KiRLxhXGmphvRHUgY+IDEAnF9BRDD2nRQFk/apWdy6801A1oSE/xbuXe8nMAVpo
jAKbznX4BG73THMyHkfGFWNKI/9rRqG6s2k8k0R9qnBC+WWhITsK+GyMXRZgpNvNh1vbzwzIZxKu
q1D/8Eecbf/uPVlRir8mXnhdtZXqRvwXHbOevrCRZnuu0DawomrTpIOLNna3w/1TuMKOTzVHcPBD
/pdHnsR5bBdtkAaYAOTWVJw4LNgSQDaClNqZ8o0fyfaea4c7/mYVBOCbnOF/CFDwyTSjLDuLwcUM
pV/kt238K4kRDg4KJAEcALE/h43q9WPtEFlQreOFNaQm/6gq8k2bzIND7TsEv3STkYegf4tZMC0b
C9xnr4+y+NN4mxQZYm5rXYFmpVn6SiLgCXXDAMzcnIgK9BcQy3ZcSbrGIH0YFA1azLHvAQ1Q1oI6
pYDtdrN4QrPo7aUSFH7dX1Rcl9g9eawqStvArM8ymblPgf9t74AoypALFrCmy2nGUM1LRLqQ8xoM
NZofIh2bhKARNVJNgNlPS/SGCiBWUwOIGdscuiMGFhWQrbycA8npjPKwOjSyPwMxeZg47pC9L+69
L2PTTzpN9iMSZ6yD1bJ3btc1Dy9ml+eO7RBqSltsMrdQZ3RyuTzsVAF7k4ZJ79wHFNBVpvFCL4lR
QKPleSwiaFQsgm/rz8DhqCFVUdKzsR/Xnx0pKXxKrTdlgLOzvoQ8XgrNs+IXL8rb6BWU2mQvBuN7
d7nDjkbAKgYjApZZ5GqkvXzFzfGeX1UGJH8JgnNpHYBQ3pjuzU1u3AvvbxR0z0arb6gVPVY+DPIV
ceRH43VWdNS6+yt1VJH2GUzIYCPepzEvRRj/QVVUy4unmjWFt1YgkQzYtuUXoSFwB1nL7yEbuDAs
R1WRSZB1heFHFkqwO1fy9LowcYUouVBfCfqEjoMQZuMUDIbDD9AgfVC6yJfmMK0awopRvudrOXlU
IJFIBRVzCC/OgsIz5tJdkXoCDdLeTIV68nfyCdI1Qt7+7Q916Z2C+B4Spoo08VN5m2Lk1V8kMHc6
iVyJvYSV2dynCuWG6R2O8FzYgpuhu5cJIbWpUgFecqKuFhN378shrfjNwM6oLHZnOReYohwXVdue
aTFDXpOFtvz6+qUJxjn6TOdjT7oZ1XVFfKhgqXHjpULh4NMXwsvIqa+zuVMIbXyMIB8QB8Dh6XTF
eZzlT0DGY9khKp7uQqsl+MhbAHzDTUy+gCIFbeBTY+dx7/Z6e0zkuEMSYslNEKKLqiI4WQBgnxob
2AUB+8JNvfMO7GGl0SnDpcwBjBaDQOKzvjxF1I66Zo/1XUNuLki5P3r2BxzVbVeE9rcOxi4+IeYt
RHEYBTvNVWsPXpyNfy8mDP+ZWcnrHhwgLs6F2JRarTNWzkYL6kbTHqyIla17GPK52Arfmh0kw0dy
mWK6rbFtRQrFIGrYh+Ij/PVemSJE4ftfVDVkDmzQafuaSLmerjH84zd6UWALiH9eJtOsyiKq9Uuj
GlDI7Esnjbez8HBNwLIVllFtOjTT5TScn1ZfXjz0FZOz9dxesndea0Yxy9fyzerMwq0u4jqo4vq8
k368mrrkzy1w4IWU+740ywEmHJumQWC8w2EaJ5JsIYk8xzjZQLVn2vWJb5TDkthyIG2wy2Nj6l17
0WuFuz6d3oVyhatmltlQwreV0bl8RZPZ5I+RN0jvgsrSKa9QpQcPWCgMhZpk92WZCPy5c0SHi164
00DySiS5imjV6lUHYT704rwnrOuzb7bQLzobHBGMGsWzr5O67D0HriLCPn5EY90vRMt8hhTuaii3
is/Vpzitu0EMkUgWHNI/Eetm7RpBEB+TF1W4PqahoAFqeW8wkIR8c1unN5YxuMBgPEBipIkebVqP
RXmsW8ncjG5iQ7/X7ohskIfawt/w6PfH2F1XJ7oFJyySjQCuWTfHTTvuCl9zedGV111S2g1NE+Jk
cGSFQVahMxGdawnQ/ytjQ3tehm2LoK0Yoauy8PjsfBFTJc1XGyrbVA13qJFSLNBcAMVnBvQ7zNaY
U2f0e+qfx8KOcc3X2QXkTKSHcPEAYrwbdY/cAlOXpB5n8MoD5hy66zgMAno/j3bKn3ROM1C/jQi1
a9KRgFONm6H9ZHF+JFBsT1X/sY3DnNsaU1N6uSiEbhAnR13gbzeQ1LlmWPzOtmM4X+KHpd0qIHaR
VU8DL1P51EwcGyedTjnAW44jsNpmf0lKrR6ySeoG7y7y0xYhsDgInf8ndSHMT1bJZtTrAdBSJaXf
rWunwNm1ulprMaCgjmIszXVCNm3sVHwbhfuFPkB/Rq+aDa8yObViiLVHkSGl3VraztO1XhJ+letG
rrjhZRjSq6xBPN+hf0M/t41kOFa/D4pzbtq/AzP9r1i3hUhOSALp21IBYUXbMfT/Uj3KtNA/LgU8
bMdp7K9HFTOrFtmC8hEl3SsdxVa0Z4q8V+z5LSne31VmT/PL4AaZqDRyLQYmcN7z1NdjkVBrjDwa
UmFLFTGVN9ZssOPOUXnoTF+HuJPAqrDUyvqD7223yMSa9eDuaKho3kH9gHEuwnmn9goQWFWuZKoC
eAEAjHvsEsYIYjURwRBJOkhx2POm586D4vLmJxk54Btp2UOvOGJpKtKmAMZnTeVP4Rf9OSTQwM8P
fGFL9OLmbHI5cmydSZR39d/Pc92XMM7P5OUW5szWxIao6PQJ3hgAPyoGwlh4pNVT/gb10gUEeI6H
5LU8UnKK/jztYzz0nVLQ34wxrRZDjcJ/1Co71EsUr0WXzltrJDxHTmCrCD2SXoivudzw391lGD3R
0f8374gfeI1NVuDuYB72pDzhmSLkz7cbElg/gaD/uOMEu9h2tr+CmqRb8fa9mmHclRQGVkgzs2ef
yS0tO2oMroJ98Zu2pRhnCAY+aSLnddrsn8MBqI7oIlGI4V+Jf27bgD1u7Du+EouZ/dxnMO/m6euC
omW4u9Y+W/PORNfVBiAnmLL/2wDY630lheB8ggGxUacg5vs249UJ682hGnML6aLu3q+lJ+e73dBh
66WstXMsWdiGtcnh4EIac6oY5Mu9PrPGe8cw0GnQJjuYnCFrCk8RIdLwxIcb8TYg6/tbUAqArXa5
gQbX66jvvTTvJ43aaiCCXJfQl4NoHA9i183Yu0pDPVAQ0Huy4iKcKFXbcZfJbCace23UQrZudD29
hKVIC2HbPrZYniUsvAqCjLezCxJbIXMt8f/89+txTJ3Kk4GiGAU92i3WuCujHua19fBmgZehItDq
QGr2eCmzCGgwFdnBPWTECk6HBJCdnOH2BaFDOkbqb4d1BMdisN/h9VBE6GpI0FVn9nY8QXdzuAqw
dBBogXaxwKkYZh8G4ppoy+HSp9FlkB+0mMSwy8BvJx2bJdmYls6Kf7maT/t/1T0Wz+rtT0PsZomK
5FvLbFcf8hkpv84/rayMzRwQ5Dr9Y4hD2wAq9BekAvj1ttrNRbXExOwrinDC2mnF51667PLccYai
oPwysEyiAZNlx87yNghmgwUrLRoqU32WPnEj41rg/kEXSkuuWInNVTZxDSBsyP27njOqfeCKbA3k
Xd7pZtPBmz/gTOQ0StUwF+LcBUZ/M4o4NtonOmuWljXTqLe66RHC12yCO6KX1a4/5j2gbwh4m23J
n7b2z/CVtZzDkNFkQD8VN3SmD9oQ4klB9ZbzdEPq4bSeZL1J+1BFvDu9s1/7JY+yG3lJKJxYTy60
WkI30QDC2teCFHyldpaVZjzHWvgXEE/0Yv22bzYddAqTYtgWsUZA1VD6CsiivEJlrHzTvvjtcZt4
f1TvNNvAhK+bF8TLA3CxaafmS8ufqRk7dAxpBDicKd6ABFNLD8CyEsWS4uCGSqdx59q+tfkdx9ld
VDWAdmzCoRKCVDugNcVSLrChYpxY46J/Hl2eTyBRYzEr/LnZL8MLtEQbxAq0Y1oEKB3iJtPjG0P5
BHiVbWEsI2uE+pBAJMcQjXUgUZkFAvPIwVF3RbKek0i6fzRqv5ciTyTSIej4XpTZ1He87W95uREo
8iZBAHK3lJZ7aMl2CxfI0YXeGnBZikRfSlHNSAEIF6mmCYQoB9jv8uZo2gcj/GSC/MygpZY9vtQl
PWqKd4go1jnUCGUU1zB8EDIj6lVI+JhaE30rZeVZdaCh0Q8ih9DgJZlSqiAE8svgJbQDa7uFOhTU
DGkzYzalkyuWwvhZif6MIVM6IOAowRowDVfgUSusn9I+fOqEG/lcR1PSfK8Tjg+cBspoMMwxeDLq
DPdzeJZEufe4tZ1HjX0E5jEBArSiQJH41+y19GMNPeQTdKyjPBu/brDb1uFfhT6Q6sAnuHXfXhyz
hiUwNPg+os2xnm/FWALj3CEe0sLk+NoK/zoP8LbOLUwrkVlXDqOPxgHLV16arxlAwLiKMYUpwxNq
KsdyFr6UodPvXcpTSkBzfBZXFNvTWyLpK89KMtK8jaMANC1IYQ6HQnJvF+xtZHCitru/eoNNFIuS
t9nh7Yb9TXtKcm5bZDYXX5HcyeHNPR18/np+JGCro8GgTxjlbhVM2tlvT+g3vOFTvrXxwNr2E8JJ
DIo1uOSY6RL7lFjxy/PkswR5oawIC7ZUvFDwrdonD1Pck60oIL5YFeacnNL5UvypKc4pJDmaogyF
K0TF2cAtVCFbi0wBaI8YvfaXlWbVqGPuMWQ4mmr7k4jI8Dv/pJvH/R3YIwftzVtPchu7mRf/2doT
oRUXN7JtJwR8URr5qJ7f/LBu82l/skJTmXnXZpEIt+7bpVjAqoiHA0rKwAxIRNOOSWqA840RTWHa
d6mz3D7ZBOq9Z5VeaC/w6r8xeASnUyQ075Mg8Owv+0tOsI+qk1cmCeuACBrNf+LHe5Ya1E9mP7Us
6Zm9yJd0Whm0cI/f2AkwRmoFsQa231sdfAB7f70pavfAi2bs2r8Jxy4dD/W30tGsB6X0hkfUB+TW
OZTUWkldg5pFB3+vkIFCwwZ5HQU32a+WN9MEvCO8atfRfFj33p2VdJR4s9jv9Ro46OPWLKL2u2D6
UzI+2at+KEtMf5mDfWXM9ZAj71M6sozRGhS7FRbId8gK4sOnfj/eLyKYqeJJ5TMQ5bQ1gHK9bhA1
lqj58absvyQkvylsmjjyqHQTGB1KkzmxnXcUSddfQmie1rFDNTeL2WoQQyX626mWlDW2aOPDz8Hp
kZ5BkvOvikFZRHvecoY5SrEXIotmAguhWGLop3oDCA92FVoDQKsGKTe1/XFaBupLRDgujtxlJl+y
NLGAoULitLSK+ZoGQ3FpqLv+y+A+mYuGJJsmVuIw4rZiGDBEc3u2VfNMwl2CQourYS0I0L3pN21X
YeBQf3Qe1X0pcOArUin9Xs1VZrbb+pQwMGWIefId7EotOeM54hp69sjf/+P2Kgl/jqiHsGoCZAYH
51qNQdb2erfJRhcg0atbpKcz2I8v6qQ/AKn/m8wPAbFfs2vWsSKACTXEcKk2SNRbh6rFvbwbRwBq
hjNUWYWtDjfLydZ7zzKY2XSX2kyqf4GbhUj8+P26YaBkAB/Ms1Dd/cU5EN1yj9khs0AepjzW1yt3
Z1gFg7OJx442t1E6KSkKeU3Q6hjBAUv6g2M7h+Y3y36EWmeIwKOY87yTKtY6Y1B2DDO8uPtUp138
oVfRMN21I9Ub52Lu6ffGzHQqM78s6KdjUdvG3ReQY9lwqexcY1/9AxKhG3Jmd1AtM5wKGp8vPLiT
lOgq8GaxUvzGxgEi5BJODxtAZsN9Y/CQSUFpTWHwIP7TiXDRL5gdRiKqDVyU2l+QY6jSdUstZbBD
v2AMwhn5ce6sae98yBJ/+2kxyZLEajGvEfDfhl94RxFn5z7zVhUnZ3/H4b83e5kZyS83adPY0vzU
RlUFePdXkpoiClK7lvTehzNG3V18OBGRIeH+hEgZOj1I/WlsvjFTDVLVu+ZemsgS0qUqxEWZOXge
op83CxEA/QnhTL/eYmFPN5z1eCkvlxRx4fc/I7AjEssvg9SgECqLtRKrzwU5Xmbd+qZeDYKARITn
cgf/EyasakgRBsZ/LRqz8oDB2omR+JxDLHzyWT5PgbXuVJB5I9C4QPDehwFmlcRHBj6JkwXnMAO0
k4tibF/29ye9gVCPWxvKP0rAsOTdXe2TqIDYj0eOaOaFuE+4ifeONvaFvORpin9zsCRDh8hnGU6G
B/HHGYEJSd1BxzdqyMK8UVNqc0k1LqDk8uxAswpeaB156cjedh2RNzkIQ697Vq+YOrVzfWRwZLbR
FK3fs5OROx16HAFdlMSW2NwVIrnZLw9ravxKsCdHMui2V2qaI7ntJrXg7CbDzESKfaABOID/8ezC
CR3p74oe0Lb18R+mroyX+f119S2Mg000ikkXchK/7hrOGBPAjxV7cUncBugqY8Q8mmmpCtYMB0zW
ZFpu3YHv4NyoiOkUT4EFia4M6xXG1nfYb7D2StDaprcN3MO4ETmzldfvP6nRey3sX7V3C2c4myE/
WqruQC/1Nw+yEEVk0VFXfrBnYNg2etr+aJlRepgDgxDGqSwc3yPNWfqbZs242z0To0+SXwHIOXsb
sRyX6pgu8qj/AvRnjvPsoSVOBfKWy9btidukgQ4BqMcN/9MpP6iT1ADPGvT56HEgj0dfW6HwCrDQ
Xj03QrUlvXa1jFQqnWSm7mwNp2OHfxhhJQTMkrWE+Cz0qlac9hi96gQH9dAavxXvkM+8sObtI6d2
8PWe9I8l0Tl+F6zCZsW6EeyXHSGo+ayuC2M+CeTCa9iLhoWE1Pi0Qoz73/WSbZKDV3tq3G8Z3b3L
Og6n5SUBC0NGja5WvPiQUBIt6LEdayrzAmEXbdyZPD8hFD0lTcFGOo2E3vpJFdNJ8d7OhuklI5Pc
IkD/uWLuy9obiZMCqETR32ob36gpI20ofDmqJ/j1m79tSVzSTvQVIcrjHHe05JJQbESiuI298Md0
S/s2KNea+gxfVQ21U0XXzkSsxX1eagv90/ZPb+q6Vq9PgXdVDFNzfzbJcLtvtLHjf4WmejqwSUIC
hAA5jQuoeCdXrR9b+D5EtJBi85J72CXp6fkK9tHBCFAaoaSMNrmgfi9j2O+Rj+37vbaeagq/5u/E
4gfMb+ppG0DVw0sOsFAZ5bCzzcLoTRbZF66C1m/tBFVqq4WGyCOxOaas/gGCmIs2cesmBBE/YbAK
ayORIj10WUCfqLnsrnCCRm9bQ/CzOrb+kc/65dC5BrIBd8BJl55uU0zHWirqMIVD8x39vZgK+SaE
C7oJ6BTfEo5zJS2dP6YfhS2cii6rea+qXw1FOkh3LwEm9Gkn1JotSCQrn2AMElm4PRzu3kYfzhMk
qzu+djU02gXko0WQBldKj7gEpIIsPaYThEH0M+B208OY+psRkJexboTTRGDYnofTF/NOIpgKxS5m
dyg4HO1Z9Og4JAuY8uBJPetcyhYqbLeOAdL+wxbLnU97qktYEewNJov8qr2IO0JUSm8SX2lNciWG
psB+B1waBN8Vlg28+ESX2leeJ7+ctPjBYNhyyUln6j0xxqv33+rA6gIF9o3I1jnYl/yJnw9dWMwD
XssV8319e4lDrfNMKeftBmAAVPwMtvzWnZn6yYzb2CS8rC3XxT0tYgFzp0rtyOMOlp0GUnKVdGcF
xIkvQWKxUAz2KRS010SWP0P8wydv8s3w0f8/qxBaLoKVMdhPubow+T+VYxxu/g4sY7/PQBK8q5gS
QLDlaEavpGr+0cUZuqx4RYTsCxe1y7mirLVl1rv55rtKDaf9XrSLNnS/iP8SBGfAprlT7h8DjyPa
wCSmrR7tmXUebBOcWePS5uZPrK2FoMiC+vV0NiVCfe0k+ehFueFkh60b7VDgm6FP3tD9e5GC+zyz
gf6lzrlBf9qm4ZthG1ob3E8/ucvOByPI8NN361XlzqS6HkoKVBYHJP4WLBE1DdJRBrZzy2YWE9qI
WbMKRc41Xqt7+JiW7AeomgSHiPYUK96t0lR15XQb7kcgwu3TsTO7Kk9pG6WrdAEKRjmxXBul/yqA
92DxlalUJps5KODAdBCEFc3YWKMrl9wPB0X/d3+VXKBCa4J2xjSRB4O2RrbA6WjHgUQLz58J0cQ7
r6XwBr3Zu5SWPheBDV6j6AXGQ+Kr1se6iqMOTD8mJX0fbdazN8zOoKfjP4x+EB2BWyMTmjsbCliS
gCH/ZqM0PmJ/emat0pYiWfn0OG3QIhGPdIUQNFAy+MLRjNLSJou6EA6WPdmk2W9g6SUJmaW7No/Y
bB4y/nBX7LUkuhwdcK2QPbAgSMAZN6Rc8uRdBAzelv9FSWz8S8L2dvM7C3aLEPIGAjpfppfGgTwN
dThiAVGpBChHS+5b2Q0wzBiELcwg0mrI5xEh7smzcePsWHw53rtOWSL0nk2cWpsf4xnxO7rinqv1
NMgxF4m8FP55GWSEZzNjqcJGxjeIZWGiDCfcagT+om5Liu7VctfqneNxzKXENx6AuZ8PBl3KYLmo
68asTMHx+KzxNNwgCzgDUGcLTLsCbshweig7dIF/BcfVOihrIMu98pKCfsRRtrWeq03zDK3HI7Vl
yv6VvZrwuKR3Jz6szxtsv3+7wLqRXt60pP+JBK8Y1sm0dl7LIGhlDbf5NbFSfBc00TzHFl56i6C0
KjHSdTCR1t4MY/iWR4S9gZPPCer3BK/At/+pzlEWCfSVE+9w5uEw5DFanI9qs7qHH9DztFzu/p+8
2/axRb71sOOFhDQcA+bFrsGHmZ8rKUqK1HLLrGtwbokarbOCdjqy7tgZmTDSsLT49UXdQcn7208k
mACBIbhE2ee1QlLaSVDH4uYd/d9G6xeFiXMEVYDV6yM+hZJlsIACotZ1+SObNJXa6cJDAqIz4so6
uKdelGaWX0wbMLecTPXaKuipZUHSZDUgTL0fT8GrPmbNIoM/jWYGDh160ZKZ/+ybkAITWD72ICYG
gQHsXMFFNLanPrvRmVivTMG/4k7mxHtWUKa9+DnxY+1P7EBage3/hIImHeIG8/BHpRgfB/xqn9MS
HSx4obJHWNAwXN5AdJIH8tpmycefG+z9fE4Qx5EvGD/D8o1HtRIfLjbueYs27jX617AoN6ABPKrz
hgBgcc1d7pRI9ax/PUbUHFWKPUHLXDBZZ6QD+XG2dLK+1ZmRshgza/OILdqNgN3NUZ0j8rmtWIZq
swW2DCmcT7d519H874kh5SCxTXLIH7gt0QKtnByrfVHCfXZSbrbTz2hcAbHBE7W8K0HMN8AA47gr
C6S8sU0ktin2JO4oaRlRrRgh5LL+iAta14Y495MZJ39jtzSCZU94tsi8bkN+Zc47KNxoA1CHCvsa
cgsx/09eVWjBT9svSHLBNHKdsFF3lFo+Sd9XU2ThlqCoV2eGm5vZnWsy7M6nzZMOtvZspiAEPG0J
/UXKiHy8MXuNYXviRFXk7Pff7gqZ/kJFEPgLtDhDwfjgCeZ7RQL8xYtIRvkS1MWd+HcBQcJtgYf5
7xlsXHe8Jm2r2TBhTe4RKBg69iaxkJBKxjElhG/6wZCoSKW6nZnZ3sABmlRu9IyxSiNbGD0I1Rym
9LwzDSXaLpfuXhvjWZtRa2xIipd7fRmD8F4/TwW8mmb8b2S4h7spjNqIOgowDs+EnwiinFdvBgIT
we8N5wcIDuyPeQdb71BOlZOGwJZK+A1rmFQa+4eCIhl2rucm/X3Nl9l6W0ZLvS6wLpbvhyX/7Got
jv477leh0j/U5TU3k5eeQdooMbbbybynu6nGsKe2Sg2K/Nl8qPZr7txuWQX69/smXnruM8tF24ww
GJQm0tKmsc7UFMH/Ss+ByHYmuhoSvB2E1zMnkDhEa4/m8lMvrjlbosNkPrAA8Mj0iPnRpewPJPKI
W2AN1+29f/9PcDd91ovbow2AuNcGs+lujlJ9eSyiQUSIcT2Jiv7gTc6Tkz4k2ehw62FMXPoPPbx3
8CTA0GF90pb/XsClSjwiZY5t7+aIDqtFc69imsHU/YD7cw/AJKIJKUgH/aPYXSiLPmi/rIN1PMSY
lvncZtLDi5OuRSJv6IfrRqiLPRqQF8lSFPDeRXHgFp2i98oCigtxSmTZVJG9nFGa7c0gPZ0ui/W2
2NEl5+0At8C5r9LtBh7D8BXpcyU8ZIa6ggxBVxNkLr644LmEEfj5CwXBb3cymoupYpcijtOFQNgU
kjVEOYOrjGrxq79HsibEjgklEyoEV5pCZsjPENhe0aByUsoiXQpXMgvlFha3cjYwMpcpr+cKa5sw
bTffOQxe5amMh7QZxHF2mSZffeE5tKHXVGX0RRYNIpmbUWOmmOECr04mg3okucAwvoap6Wxhnf6z
bXwmri/x1tBCrOrlNwrXRK8aubu8iohEdYrC8Iz8K6FsYPMVp7BRPYOEBO0xA6oJhKAINt0XiAD5
DXsNPLAE/8vhdGV/uULJ4Q1jPFAfV+IH/RSc28R9YzO+h/ICQGa72RNjnkRjuv59rkGG3wWAVdVM
JBG4J9u2nye0ZGa66zY/VtMrkru8tFH1awoJXUCui7dmSYe0xXrHG0ceEKCmQ+uyFEDhGX+mHwmY
V61Rw4IzxMLM4XLyJ8QUKCxAQWGiPNh1Xv9Oj/oXwHmONNWnd5HMsMQpEmh2aISy++NRVvYy0o5r
jPYCnt+MvpD/0qZNWzS/KKQ8cNEqc5bgI5s/Dh92XBPpC+1aVs/OzOyFEnglbziitRcKEPgp7B9F
qya/JifL2/LZmAxsRjNTKLW8P+PgAWmsDJBNklCYfNZUpbMw5Y+qbSM7YV3jWGZ1c5p2gtQDu7rN
D6QBNpNzq28knH6xB7miFFGmbeg5NX6uL0W/PCpOaj/TQcKOWhTsXkeoLUF5+PDrDLXpwJ5J8Rh4
bODYYiZVlFE7jUD65/jOnAev/sk5Qf6o7Utx92j4FLjtoJQR48QuNlLzjnN7bMs4yZ3EeCpwGxJq
89EeftKjDzo3/AOMNl+UoTNDOrdXCKf4/DKZTgGumrIIwCttJiOKSkIfFf0wnrMvKDwRL4ZekhPT
AOXadjQBSIlLxjVM9T+UNNO3BlsdrDOloCR9Hm+mixkU98T7Rzsrs8aGOXIXkta7IYBGL3yAAC5w
EM++d1t6nQJhsRD17aKKeEOqaqaDGXRhjludMcbRIGQ6K5cp72rXsX2Hr0mz3gjf5u7fE3uJ8WkK
2O97mj5FBs+yJbN44lzZW9hN3uK8F4Hk4WQ7Tbh+iOfXkB5ZfSNeFeVFSXa78KhlknqdXBexcvyW
IpIIcoaFiEDtGwwSv1BdzcFp34fp41GJIrXyZnDmfa+tcyLsWhTHhEFTxO9Rolls7jeKMXlRMKzr
YOG4TahMJIOJxVEAeObstXVlIzrTt5/VgaxyfzqfXGXXoBArHcpZwDeORs5rE6CwZdHL3fhPcK5C
NEDgeJqyyvWs3Y7xgt5kqdlTwIpoRf3q1zEv3viYkKZRZAFDIKPHts4F0r9REQqNGUo+Z0SthlKZ
8pSt8JFil0En9qXfyhp7Q64oTnDUaXWuV8tnAR8cm8pRUt8tyUf2UCyVoOzVddrRbs+Dah+ocwVp
yLkWFSMgH5LLwoh0RMba1u7wSgGuXB5ydOkb5JeicDLFUW4EFVBs5DvY8dFhVelBpLrRdEtnww3x
5HIEviqIDl8dp1wh5EjhN0PAcYClMPn1DOly15yzY7sJN8DGIFcgwBQNJAy0p2GNtMzHWYUO7hzO
/XYgjSHAf3yJs6Z92c1CAYBgHS3OmHcOtexdeM7rjN3uhpF6BJrKSNLgHLu3GtiHTmzgK3BtJJEe
tDcsSDMBqRuw0CbBvFubub97+9vN7HLIFSI1jsRn0p2tjy1w1zR/ZZee312aSNIzJcWmDpN1Yd8W
q2ZHW4QS15ASLVDmGMckrwHb3UzCYLGqZSzY68tKKU98xRnI3JuuU/Ifo9GWEvui7uZc5JAsMFzv
LKymOawgmp1K9mTncvFFc6Pqk86HenmOTf3EhSUw9pPo6twXCXT5S2kokTQFpOJvdnNQd5BeGjCH
WmIMwCLER/Ym1nDC/FYko6HYZCLQOiFYl1OOz9/f4tafU5uLjSiSYrVR2c2OixhMNJCVkVgZzRiX
9r6hIKY3XXHy5lNMgj5wlvgZKbkWhe544f2jXIjYUPrZqVEyeHAwr3E1+5tzZkfy3Cmmn9QuiDsI
EmZtg/iXlSEkYMVR0lvylJXZUEEwtdHLBnPCQPCCNWlUA22e95TRHViL4XPUzu6jvsFXEwvDKsKH
0raPGzugBrsMghY8BGhZ6h2cOfqjnQV1bOHZppOPbLkmrtLDYx9nOkH4gH/TYLEOR+UAHy4XvJgo
Tud6P8FlRCjhhVMImdH+Nq34IFd0QU65SFkvTKrcfDNeOJ+iXAHMbLCUBLSTsFl3o5PUd53TnkSe
IuvTQUZiAkN2WivUqeqx5wghan9zM5Xlg7/uIsZm+L+PmF012pS5pupEGTaEjqoRHrYqNzOS2Iqa
/nygvX2SJBnqJZpwzpeaDfJMZB5MKo6G1SfCfg5QXAzww0Vma3aXvEZJwwuOvWPHl6a3UWf/dmTC
3v7SFUWUzAxqe7WgrUXuhE2pLzwQQowRjesqcYx9SvoaejXOKlFfxO/cnRAyEuadK/16PBHCHw5d
/hAZcT3xkJdKEqeF1AdEwaj3SUyil888zh6z21H69V5Rpg8N5ixx22StFvdh/730XtPDP6z4W3uP
LW+fTUGTySRWh4qNN6k2+rDf6tGjrP6yFBQqE8hY+L+NaRggH8l6PEUOTow2JfGPP8AYyyDOylUM
vICw9X1U/cvPjLpF6Trx/FKMrPX6He+b4G8lzZW0l4Cyjgk4hTUgoiUIATJFZPKYXR1vbf6o4Ike
7EHpVnWuRqCcKpedf77QtwLH6OI7qCsMaerDxWuu2o59dAcrr6y2hcgPZ+Dfe6OJC3Y1fxe598vf
a7vK3/J/V5HsWze6T5ixgNX6fcrQKeQCpWM6oSVqZG0LIiLcUxEUS4ozrAxn/icsTHGxC68HOwkO
ZJclrhCqslecUvtZFjRNiVhJfqYjAnrE7Pb6c3yHgMgWRg/YezIFtKCUMAq4YZNs1wVLng2ajgGD
nDRKCaPa/FdQQGGmW5DAs3n+6Cyvr1ktNfUbRKKs751+qWJTAGJPqLFqoDw4p/HE20D88sCOZih+
BgP0XQAFc8NwtogEoqOMNd5XiM1x0AZu/hvE0Yz8KraAijgrGRrWBqtSxGHiypbpBcMS24yRfeGU
HJvHqZtVU0Jio2iQV8jsErJJDIoNOEAfx/plfySUSB2biCDnddy7hDRwLCqlJNOiaO3tKLr+Onxo
aGroMniPqaHFotwqY4luNEmaEeGFH1ck2hA3nujUw4T55Xcs33ET0ypMpyBCpIOhoknc9fylHZ8y
t22LY9nxAuc6dMgBUnwsDn7zZ7nvmWx9DuqNgw+HAmbqDTpmiTIIOkDIuoohuq9MAr+DeInkdwiD
39MxpvQGx9Ci5vTNgiBc8YR3//lQA6P5V3j9mA/UR0jCj9nX0cT3hpYVqVXNv37cPlHe62zHFlz3
9yIOLXt7Sx1u3/7l2wE+zNsQggPqe/gLGvtGxo29YEbyOuTYb2dmiTG77/moHkfWKuczcSrPof0/
RxwyijVmeGpOHWicKUWmwvphKKdUh8SfHjkR9XJJDVrbShrcLfoVi4+7NfIu7Ptn1DOpNxQtG06X
EfKo1BeEDXwlFVPCqzuvL0x26fzrMn8M8ZNqaqLOQJEKrTXX2abvjKFV03liinBKcvL5I3ZMf7sU
B//eDr0mJPR4zM0uOL1rQ3ej4M0YjsRokNyogpYl5eVj8zie7x1zNnxbiBLlupaPhf6n10OTv/3E
sLQGXiR501VkEdLz6/7TFL8elTr+FXriCttUkRMXhUz9GX6ANpYBg5HG3ivuhKO7CvL1js+GnM/K
Wm3EopVpAdqJpb+3zSTYwp4uxDTleMD1RY1TVczWBlAoqJB5j3aTKKf8uk1aTh+2uzUYSLGMP8sV
jhPyxdKZ1dq7mGPEl8BVhIMmtErWWh6AZ8OqX829oBilmcoJA9MqhEBj2e87AIGyPXgp2MZ7hDmE
+mTlwZp99BRjH3/kS/tvY/IMWwbqQ9iXwtMs+0QwjeZa9ClvXdSA0QQn7nQ4g0DxIfCDqeOYKtKP
DK4yVHeVnkzikluQNu2JFKPmB7CemUhdyw5V1Sts0l8zmN4Y1dZHGV9PeczO3dnJ3x3PaMha6E26
loZmQcLvrxCpaGomNgkhp4eGG9pEB8KwNeodzzjxds1okaFhpJ5kTXwmOvJ8DaUEI0Mj4QmFAJVX
SldGtczD1J0stCcZOMpoIlfx6GRKguBf0vvwPPxTlVMa/EXV8Uki8HTGMAoM8gKGeXCuQ0WXoW2l
0HTJKbMCmhWMSeGQIPslR5lGKYOFEDAipMv18xqytiE8YsWiilZSp8Z4rAOsTtXPiUaVv0tDxxIN
owVF74p8fW1wWRrk2bZIqLpbNxMXHLEBnsmLAg6O7kppeBmH3Nx4ijB/XP8uX9V9fbOn6GU1SjeW
RlmehruF0j1Yj2B3DAlAXFNoJeqziJpspSsXilgV+3pyJ+WWNmO71eaMH5c8+ehPKY3/2oNbmuOk
ltE/zb6sdzIJDyd1HVUgafVLhMRwzlRX/3TRzNpFySPeqPBKEA1O0AYtF+9R9sK0RFKH7d5O2WWQ
TmFEh4D1wTUl52ko0Qm1LfC49mV6YhvNlRt4AYez+vES6G8dcgv65gpeKSJaSgin9AHyijo5RtGK
hW786jVOPhNumKtq6ZLYKBkqM4r9sgk0qxIciWhfFUuouoBFhf5AMwgeM0v5o1kEDUaib6wcza6r
8tg4pZV4OoySh6X0MTi+Kec9189vJdNej0MAG63UOC21RZBkBOStUvvEgCM7N+noF0Hedm/Q+CFQ
Uor1ezrAzJDdH+hlNrJnm6X7BuloQRWCFR3cnvkoZ2yhXXf/D55/KG4dtyAlrW3EKz49vPhurxsL
FtLxQ/9mVbe7Da3z8uWNl+OUUPNh9nnakjsMk8kGHWQPg/Xj6Fz8US9LN+H0WAMARMTRHK1Eaqu2
lvF7OM7n7ct47w/q8LgGmvRBb7YSZopmzU05vOUouDx0a3H398b7HV9sFaG2JZIwo8vKT/Z3tppe
+63I8zynwOkEjEKN+XQFlShTy2wJi4W23OQYcsWFek1+xBdqOxgIKHSRxZG+yPq7E2Ju5sDMewx8
Umw3pOCEHUSwaL2jn4p4esWOVJ/9bSmD7ppFBRJGak4KYFOJB9+M+Q76LV6P5OLX8BIJZFB7sWVp
312bImEyjGS/ZI4RR3C5r85zrMO/Ovu0cE1jbyY1H3BX/xQr7YLIvGfVl4B6/2vcVBR1zkFfrwi2
ei6VHQa8dsxHiNkYdAWniWuf9uREl+301bd7pm4av/1/qGXXFd/D1WOKT4ktS7bKYItnHMCrvKDz
9KhiZcsEFQuAyIT2V8lfOfaEDNVw94SBL020CbPm9+MwLWKYZdQQC3Tg9RU6Id4riiQ5D4IGxCwR
+vreiUNaBKFp0U4/diYJWeYZvuCyoRrV0PX2JzRLH/ghK+dgWH7dPd1AW/k8/RW9Ejso8dQ7+Doe
Q+YuUQC3FK5CjlOvrkzkxtNqKrcya5+ah/zLwr0hDUGnKxbmcoXerdm5/1lJzIg7M5F1QcDBVf60
8yWMzyxTeKdbdH35AUvI6F8xNqOTjOimsTuu23rveEG+1B6ExAkPZAAgW9VTI+Q7eDiY3XuNGO5t
zkgOHUrKN3zUGQko2aEKEI8fPjyS22ouWpPV44tJ1uI6KVEigFyU6tgKUhHoytHVtKYL3kYN8TyI
ttsXDLGg4gL/tBLzIDVXyoEUZHpYNztoFVQe3N7hWKPIooRMZMakPPBRukBmUuu/UKZ4llsNO6w2
YM+wXrfVfEJizpDZx3vT/Byna7o8+iVW8MtaCMHM9e2PtEDHrfxbGfLsl30dT6eQTDT1AD4VuZ8L
syRtSiM6ZekbA+S7a4ANXynNO6elko9tTFYpwTmWOD6SrYacDWrhpRZjmNIq4qeEPeBSD5ZK5+IT
hhIRxV7qm1Hp/+RiOha597xqLv6x3aYNpZLb8WldlVo7tHw4bjoNpgqiz08PqEvVD9+bdxcok4mY
sDnNiJaeeoI5ITSRmfZPehp11Hi40GsC9d38d7uJCRW8o9VUQKktMRlWCAAhWA2kAw6b4+hI/Hqm
tP7nld8Si/uBhmX2i2MHMSFdQgTiUghMnhiKu/5G+sqW4RSH2che/1brBqlcm7f387sFCfqOLacO
J3lepn1VJUuZzsapI76d894VBJn0K7+gqQUKcXWpUfRf344bxgxFyHLzja0ZnFv1jUQ8GT+1iisq
XjFH3RAt/o6hJGCiCBele+V3T3y91qdTIZUrep5NEF8AljjRzikRTKS4Pre0EviNViHxN3Jp2KGt
OYRiV3ARYLbWmxM3CFo3geojGMtZZ8t6Yz9sycz/kUWGiQkXK450M0jFvDMX5pOE/o26+sgQ56/b
bo5qy76eCXa9Bxt7zSIIxPhCMWtM0vdfqK9GHUBJJKiON7izyrJa4OPW/9+14P4R2FEhzKoEI9HW
Bp9gv5Rd6ZTJtRmDvoMLV1/O2Pr9T61XMJwzLE62d0bNVkBlzqEedXh/6gjcXPnRgGBFAjH3ASzU
EDy6x3y6DCQJuiflPmXUhOC0X4ccE8Ogplw3eoYK0oHzAYqPp1zOnGlGlIWegfyoolgjmKNGbvTD
3rUwROZiNmvYa8mBgk2ksAkQHxEievq0pDfC+Llye+IqnWx5aaHqUbQgdIq0yBmyjDqmvUiaFK4g
FiMAs3V2Z2XEx0aet4MlIPsA5+zMjv5H0wUAgXcFC1Pga7+kY/OOMabvIt2G6SNmP/CV5vrlq0LY
dTThXfv9HpmmXNqllQz7ArizgFQT9Jnoqs5YvHnBT9ArDuzu3Y45H/+a3XaNcccyhm8iHnXwSOc1
NkJN6kzTXAe0Np0VwOaxtnnO64zMSqvi7k6lsXbFYynoAAxLIEHk8ahD0hA7606UDuylIEqceowj
kjq3R8NHa2Jm0xVKLl10oHOjQ+b+D6lzyeN/5gTOur33O4bQlWjBGeHjWOCxpiH1JU/CjQwuuEmK
JFFk7n1NOY34by0pq9OFb2R7JfNK0TpOsW+Y6vdOlXzfLb80QjcNFsJL4Bs/MV5VfC2lL1wm0tz8
FUFkVrDAx3Nl42NpiO3q84G1XZ0djtVJTW6XS1dK4YhvS+Gk4+teOFI2s2eDeyzN8flOrHsw0Pda
L3Vvuq6nTO8WHxWTMXpFqq83ehGm+D58SZW+iAl1C/it74lsm7n98JrHfRIBg27K+TozhgUFDvdE
sq6ChWc1skWF6j5GY8yBrOMPePwyTUhLDe+eztcwT518WIhSsjjUq5pyTRBgHSGmCAISrztKKLbS
Xn9i1QcMH4GYCX3z/YcPtSe10DsK2cy9wWv3nzj3DB3cqDdJtujA9154ZtRWJAkR4vBEOzpkiQ0r
ulIPKu58r5aS0tjglooKqm/6OeEgvZIHxr2Cgg2PukBDlW/JqE4iL192qSyeRY4oJpFmaPqYkfJp
08bIBsq3/ViJIuNCoMox4ujgUNybUSUQY1sR24O8GD+9EOUWVvytrvEfp4yKB7BC5/WB66myn9G4
sIoJdqXp4xb9D7SiQ/nHuyc3lhsoUmLrkcLAnaEydHDx42VIBnnJylQdO6Wpc84YWM9+XJjYCMui
dHOLf33JhaAOXGLXWl3+D5uWoRCM4EkcMWo3lcm2p9CGHgFs92JxuE22cFjFslDVfMLb7Qcy2sh0
Uo6N542Ki6gY6eUopTNVJCxGh21HEdN4kuYZn4yAKTO5myOfU8pA0hDe83vtLq0moUvwSKSp/5dm
jXZlNTIMELBzmGB1p3CA8xKPbvIh0xswzBA70Qk/keOaHE7/cG9m8rfcGSoy5o9x8DruggCd9eU2
T596AOZSprz52FFL1fm5BWrhshIpV+yjvVxDvLxk4yT7o3bRNnLJScLH1ifjLOTtxiB43UhCLIgB
QfG3xMPBUVhyaNFitaBAdPn7YfEt/0WGsZ6W7A8cjGTn5zd7xW/Ro8XNbp85h0t92Mwsdnfm8dEw
GXKGlaET4g3gtpoGaFd11DCHE8ZmsQ/r+c1+zFp2nDLlPIV/qffaBnV+Wl0PX9nE5B7/mzTHuElO
wAoFct8R2v4kbf3NwHRro0C0YNPXt46V4wiUYB1+I+wjum6QfmZQJXVj50ezyjKaWmCY9bT8zv9Y
fXahN6j+zI3yS5/YdGg7K7xU46qOMaoCSVwUBxMosqp+KV4QLWPaviEfNpbYDavMNiIWBUFK4EzJ
CCsIaSf4xkDlK66NIxzT46DIjypa9Hno3tW/DGqh02QyEQy/Saksc3WVBVINkoO1xIqzi1os4xYY
PLe9GhurvNNS+0qg3lCLgXfzBKWnObsDgq5b5iyaGd7KnuX6cOMIXI8ACxM0Ha+63HdXzykgJJRY
OjHjz/lKBTIMzhiCyVcu9Z0LUJFxfl/LsnRhDLiAsaXXNNHL67ZEnTyDuvf8IopnpUjOXYQB9gTp
VZFGkSd9pvi/cJRtwEscJTl5Hx3X9Myc77ReL22omBeSuaAdilQ/+jA1ZWjBq1oVoWuxydYScjuo
a0TMlvI28NB2wccjCyeCzQqqOluvFFPfJo1oBFDyu8rfak4cYiPnwUJEhpRztQsP2ESbz0aCSO9N
GurGNZMgyw1y3VoGBCmuBInVTCHzZQTML4N1LY10Xq026qZ8d5yjxMayqRE1lmDMGtK45lIMjART
t7LOB3fRgUKQsNGvp94QotTuMbisqrgIy9/w02DvVG1g4VL+QKOmmIFVwlckpcyHXYKeAl3csZkW
VID5L0o6Z7Vzps4MdnYOH9uYV4b8MCAxwTG/omROTrjvRhCf05IsiSm93lStCt3EFQp49V5ZNBH4
Iu1TXDWSp5P24MRxx2mOS5+i7aBhdw1051JjZ2hYtMuoS2KUvU1KngU/f7IIu7ljH2tLXg86U/Dh
D48vF+Dv0ARE+5pynvUhGsw8iAWpnSA2E3gpqRSzqlLKKVOv9l2W1ED55foa+kBXSlLj+RnWp0/o
SVek+o3H0y3yottOIaNJK9t99LfRuOPB06hn3b7BVEsy6xEFqGiA3GS7BIPirJxsId8GMuwGmxkv
HsSjQZou9TMQVJ2vj62nVSTgwsdmJ+RVbVhYq0m3jaCLVrXbSF+htPl8g3fJl4nUTV2FPlkvxq3q
HNCrEesk9JTtVAWSJpYXLz86tK2j3LuUOBew/kg3I5n0ODdFe9Ur5Ud8rRPLpnCGfN0Uv3EN5kHY
6nL7o9uUdrA+197eoOcFeca3fcc5YYtw/E7jXEkJJ+VyfDlh9Na0z11yvhLhNdWUZBMa6iqGPau2
uYyUEvWNuWsolGOhJJuyYRUBhlI54YhA4OqNLnMPJEzayIbXLe4BNql/Jf4/46p4oX/pxqeZeZfT
6ORPid9k+6MkpCLVcjJBWvCw2t5RJXRJHhfqQcFQXtcrPlts72LEF53tIx+HMJKr1/t0Ahdflf89
+JaDuEK7C0L+CBaD9HyW9iA0ogKoBF5fzIDpXqNYLTBvuQnyKsb8BjAGPJ3116uBDGEsJEeu+/rd
oactrm3FnjVrBzFZWAE4HRk7RypS+iROBO9I252CsdF/n6xgvGKn1vo7g5enalksLOOqsemihgsY
M86lCpqD/rQgFnVkU4XXmsAN8HjZovxc1ShUiMT5FRZvfhfoTP3aAgQzXreBc57bgTxvkyjO/2T5
mRqnMR+OGrilojg9poM1vZP0lfhknVqPRkb/w35KEXfsnZB4yB29urXnIgqDZT8+Wi8PAfwhUqwQ
ExTelm5ZJk5H/gLh1l8YjKXdm0jPUW/gD6JC3cuwK7uqfSZbGEqljixCBHwYqUlsWHRvXTyfIY0w
6OoGw5lVB921uqZwsbZQMOHykQW7yDDBpF+/gavAYBLUa07/9P932lTsmQ9ZTuCQEdhiUZEEkKV7
jAfr2eBf8x8UCTQkCS8sKgmC7IMoMMtsP/56FhMfyscV/YvsL5z0XGkw2VUdyBOZ7UAInAPVv+gd
W/zJG0qvq1vW7PtAqWe4Prehcb1lVILMibpL7jmNDI6uDWTm4fVDBPJjVewiwonfq43T1STukBJa
q4idpM4M+8yb/dgAs+6NgJacF+2e2qQDQ+LU6bmFsyn8qau1IWFgVVSk8l1DYc9OlRimpGKGdrf9
MO5KvSZnGqaaIDnEoPVNHP3VeKJJjgRL7qzhnIGVUs3tt+jNhz15iFcpbmECUVlMfKxWLwyn4udk
U8Vrtn74uPCqHs4pDuhaafE3i+JoKkOPE1KHZhf8PKThlFw51mIyMzhTwrYqr4a+l0tRmtVyWZHG
UblSPgFIWY45PW3ehF+Fh4Y6MR1QajNz9xLa41Vva5li5o+So59r40iYM+Z1ftd6Yr8/e4TXncGD
clMBonjv5pGiXdfaKq6/8gva0ZI+VKD6fqA+AeOXsHu/uIattkrYwkstzCh9AQXiAK1psPFCR3j2
5pZucPZtMWbUxhDss2xfZkoJs4xdIWLt9QBSws7aqjvH90umHJIEjHKj6rMseS9fs6EBz8lbmmVe
flcqP1+B0IjyAtCDbFTZUBzJYxoM6t20FmJGcV3ji7VshHGMZRMObr966gyR/bVRGQ5DFIlIgk0C
VL7Ee7YU6gJlr5XluBuWMs8FKFcq1Y9wysU/qglKOXCVjanMOXkc9vSgyxdfv6Mnhg4IdMxiwAUJ
tnI1PYU09vs74kJWmTByaiW1f21DNiTwqlUgJ90pOCT7wWCpTJOBsZXTLGTrVxIMW+tQOWdf6i3y
/vmAM0vxMXdQIXPGAfCqxGZWWRtJDIhOywAGGJKuylirKVpJSTitm1OEsiw6ji8cyvFYXRhHKqrM
NYDxvwvXmIQUIDKt0Yn9e8IEBSSo993aRBG19bioJBjatr50lQcQwdEzi1OKWu6z85jbCmrdcQ2M
qBBlDjCmTqCX4TjdP9QjTera23WhqB9aFwjWBAz0t2rbzkPsXFssdq0TXUS1ZV3HipLK+Ff5Hx52
RsnNzoM+7T0FUybQ0hfVpelNzeU6/iFj+rUW93vyWMTSPmB335zAgxclmjGkV+7yRr3sRyQFe/lT
fZiocV6t+YvqC9yi7iHm+Z9+40vW+P5NLUvIAYTsvS6JXfxCj08Y26IEHRCaMa7Uxz9bagT8bYio
1vaEYDmCAG0h4994emkybmKTFWWDJROR/2ocuKX4i8nJXKjNdO0sDhPshhjmOXv3bT8AYmXs1eLP
gwowJKWu+FByWdA0ay15cfJofh2F0LGbCIreZTNXM9iwYoI3En8V5Cy36J0d0emrno7xB0H3dzaK
c+U8EXO8CUaF3mrf0GHTo/Hcd4DSK0YpX/yk2ZmIu6vg6pBuvBnFcGcmLrTvVRawwWs1GP1UzhyG
dplxbunK/lBVj9se1cdawlMV/+qem2eGpAIche33cPVvCNXi5x/9ytI78yE4wRnrWJfa8SJjjfWt
eV1dD9lId66Ag4Tgxkri9b/02oHZ9taulvkCYWuDcI+0YbR4hj5H6KJjLsrjzx0IwtUml9RfgZ0r
qifCJfQD051T5DkxJfKBlXoa7ogSg9ZPfS8+YvdiwOpHg6kYTUkpuVN1GUCD0C/3jiENxqvDe90S
QzS/8p2r2XHSIRlVlcIWRBTDg4Oz7d36YxDO+yp7SVGANF1MXhCfQyfkabUzapsdQK6V8Oq6Ak/D
5dKtsi1NCntdDQxm1aHbSbnPJreP9m/MisMZLVGEAMV58+tBdF+vvwUfU2D9q8X9h8QCqxeaQWCl
DiGDs/qHRNAIu3lub4XD2R5rlqY09F34wI2iIcmJXZfMV9MawH/2b2WYIJl6VWwD1E6KVOlvK0tP
Wm8ntY1/hlfxJJuswjXN7CzD0MDEMYKJYxpuNgvNK4uLV6EZapU0nYCSsSaxQBj0Cwe4z4kDdsbb
eH/NmV0fOvTOUT5on7WdNXkjS+34mwOOpGQ35aoB5LvwZsa8UMmXpF2KkC1FjhDNGgr4YdPiwJ77
MQDIJCzOgumVLB1r3BHj++PmCLQ/H2sW6OJrDTI0cYbviktfY/X/lJuCcRzR+Uz94VMh4/mkTlJ0
pB4Og6h24DVzjDH1a+S+Iigp/nlxu2Ohz8iAIZGoI+FbkGLY27s8N2MicmlOhg0WdiTy9NVRwGeS
gcmYmlIRH9veKjVPMqd/Ci2w1DvqizRD+iYn5ZlOi/y1JnuTCKCtQOJaUt0/4SqYshW12dvQ4NSb
MWw9VN3/s4ogPS0FoIfqEso6LranYCQPKOTaay+A0DRQiR8lVxIuuyleHeVuJTaVbW9VQ7jG0zf3
ZX4z8aCId4YPXqyoQHHEPoQYN0RrO42+3uJPLppD7OVv1Cb+q96hJb6RZu47tEF/xl/4PpzIQmTk
LLnYV3GJnVrdYmpFGWZMlxJgmoA2Dzm6qzOir3+czk8ziiQ76ZMoLdr3egRgn18H+xxKdAqA1BiO
bEVmpXLCOCC8R2qX8vZpedMh2tpURhyDDri81TDAVtA93qhV2b3+OLBbFMVumpm/fnqusfaONg7B
37rAQkLz+W8b7DoOvzu4vk6cenTnC9EiWPKx5CqFVoClTfavmXpDWjS4zJUYE0esYAiTP4Lv9n6S
6YnQ5BL1fkIWOCHWeNFjQqeFKYbtCjUhXYXNn3oF7PFKK0IZ3NZEiKFoCE6Kj37r7ZFcbOpYt0ha
8PlD1vvJTE/eoJPmo0xIXWYHifj4a2rmPu4SUoQcH4c9/+92rwllRWMjj/Re7po+vbeuDHsY3O2G
fCcxvMLPLv3kE7ttWRLYg4cUNDgjBNEMDQ1a6GNNv68+w9hzWN4odpRSFIJcG6DvHyhM+jDdbuXR
ZEPDBDjBoCYSpmzPDtLBSQ0ItujbVQXyMogfr7qpZXfHq7MwpK3wGLwSutos0IYpq91mZNDawlqF
xHblAq1HSoxbIa45g61oicYeQ14hCojxI/iCAFc/B3EaG24RyE8s9vUOPbwxUPHGYpHGsNMP5Qsy
V8efR3dG4FemysfcuMk83W4RLSiuK74ifO9OVKsrMl/EdPoujbzUnuViEIgbL3Zkx3Jj8/6Mt1At
YMo4806QBZ8xDd2pzm//4i4PTdXKfAifH3J78gyOEwL+awvutqEDe6WYMBZMzR3iPSpCqLQrj9Wp
P0y8e2MKVqQbsq/T/gjy1rFEKUYookEo/jCuyoP/WC7LLt4weMjwvccAYuaTR3+LR/2/X09fNSQQ
EIgZXlqH11bPogVZKYtz15v4KCSgyEws43W06lmHdOtQzAw7LTLsGve3UOu2fG3JzSs/IoxQbpKU
/r0VhzxRL8/5n5aFTg0Fn06sFeY3xOAFEk69K5frTGX4e/EpvihFoRXwwsl/dLPTAp1zA4rc/SIP
RjnspBK4gtGHltKdWBCV6r2v+kwkOAK4pkyf/KJWNCZ1YUV0r+HzmwA0rpLBYWUFMTlJdrGRhOyy
aaOw8sN7JCrBc1UTewK/1Zkw1lZ8TKGNNZ1U2PzkZtpEDDOJr/h0/uf/HSTZnz0D5WBWYwT7lBxL
hszxMbQhD+Zv2nENvY/Fuds6KjAW9i21BmuvF1Rqjpcy4jq/dxSaWq13aMr9KbUpCkVCP2iahvUN
JpefG8nXsepO0wBr5NT6rpqXg1cSPVgptYUslrE8KDmoE4ucKEgvBdBoBTCZbwHlu4BTXLI7GLus
E8VXgusZAQ8GBpgKghmC5te16mxDL874TyDKnloB5HeUi3iXHgQOpTel3T/4KEvUuV2GujoYIU8Z
TASPcO9xiEDs4klGBjUffwjO4svKbZTyOXajhJiEWgAa48jYCohMM6XZOHrcsYmAfctZt8/7OPzU
YxHH6YdVtFpF7zRx4NlDZICgxwuntp5Z4FmyYMJLOZr11BNb2Bxnrwzo973BWaQ6/eSNpqiq29fP
x3XTU6yZtjujU7QG65BWWcXl3e3F3V0LDrr2flQ/Ew3Tr1b//X8ie+nCAnKYshzavWfP6fV32SOn
1PepPI1DWy4OHgKaUk8/vQ+jREQ3sAuu9CV11BDCmt0EpawWn+OW6JNFuExkaJ2sCcxBlX/l1Xep
eKIY4FWLXezlqP/H3aCW9abfPjmXM7hqtKc/DgzEVaEkCAxqd78Fa83ncsYZwr3BNLNC9WcmlMI0
UModZh/edVikZWcAyWR0ps+j3fTU6D5fV+dFN2KnJfTtz+1cMD7+5foEOZq1NZUBN0selYiYj5MN
3NKYqT+TYtnHpZzUvqTskASo4SwsQk5cyPnMn6jgtDKgeXPl7AHT4KpJYGYizuMkVja50uhSjlJm
51da0XkXWSCW6Is5yg4lEDUUz1fQCpjOVXltc3lCoZq+sdHrY08X8yIIxtDgafV3aZw2ptJh4/kP
lp8betaiYQaARFEWSSb/AGLPtqTCoPI7Eeh+c4rZGlScFNo3QZoNlJ9yCBweIdyhDvcktTsNVDWc
BWigpfPY+UUwOgw0oKZG/7uEk6H7Ukv73YltlXjIy1DO43N1iRYApsdAIi2eej5QxSePhkaTVQhP
u4tZGHTqbb8gy8fvYoSw3s/i9aXE/bhmbY3elcl7VBhi/Vp6I7l/bvCyJp5I9V8iyEreuE57kf3d
8y4+jnqTS/QfZE+FAcActoAg8xURnf9OKFO+ofNDXJslc6C4s4rmebGaQXemhp4P88JMmPEdxPjr
F9/mLNWF/ABumiv8q0T578DC8cSTJX7z6ebVYBveE2HKvxYojZj1+0h7o+HH/59Clbg/rnBiaaCj
3mY/GdptNKXfqIHtUWTuFiPyIocgJ9vm6Vrnp57uCX3C3CUH5axTufq+Vy+Lqj+dth2klAhav119
XIC5ikqkvCsgM7wukBufjmnsGItS08un6PBEmzWlbzhvEGb0/qI1gDpZj3Bo73pUsJaDsdS4K8ot
kdMfMBPfSGztoAws5dKewvWjXmVZlDMGYNiR//iw33lbAQRNGZi+PSIIkqAk9RB5SIaV+VCH92vo
zaJioJgq/DlWnE+Ur7Hd7ht+MzdEIcVaLfCnvIjIKD6RaQw3JxN6yOH/7rJJbQDla4rlV0cvlAwl
6Iqid21XNnt1KpuJoxHUhfB2TgFs7AHvkoqqQawDPWLR09ok3kZYeThbRZ2kvxcP7LzWnN7ArkgK
hiivFq77zVm2sI4ZIDvBsdGXkaH78eV41P+CyVgHKgQybW1k1F6jWI6Fb9tMxxlRc/OwoiIw0UMC
SeRbD3bBpzR0cDjwBewa6t87ffxaRuWfjyUN7We56q6l0rs+NcsLR6/1ulCGGjS/midmH7dveAp3
Z/CMg95UUBMrsuAwu14oVFqmpPFOpimhWmM+AC2ZQu+Vdvqfy0KxIZ2Sp8egpzupz75IMNGJ9Gsl
Kj9PPLzAQaJL8SBhy18klRQdKJmNN9D7AnmtRdR+vfB+LRkWJBQvyS24D79yUDY8PD2wCBeOLEzw
liX9JiVfabo1HrVLVzPjA9kq3ZfN+ryfKLo7KLnVmND2NNHJpPGcDWBDDfG/2YO4LYLd2RL8ch0n
JT5xD8wPTebdv01AxTdFYjtUpuGd4dLGLE/HpPAX5b0VWT6tYRhLydekeLAhy194if65zbjHxc31
U1fC/BtlQ72KaSvHeKSyAkNP2IVm+uno3d+66ajh3wmC+dGw4FuZTf68qgR4y55mbHYpRxP5pgKz
rOV165I9z1s6RZo4cRUehkaMtQadn3GD/iTc/JdM/6gGb2TolZMU8iOassCIJwkpfR5yv60z4xhh
q7HLoL/ivPurMfMaR92aUSueu8rUBWpmZAch9klKOtyd03kTCxQQqJUvsfGqcSJM7qMkVE+zvOh8
SVTwiVMWaARJxAXy+nrz0PTZ6LIp07YdoLrczcMgMa0dkHwCbhTiTotA4wsvMe9Eg/SV0IorIIoF
+jP8YwhAcWxPGHBsKhbgoq2ZqBGNQVnJtgzXwgC4Cbwp9As7LF4tVBPJqh7ZrfIALpkUttx0HDf0
fcg7LF/8QdnanEi2Cxw/3HS+TZG+pi45xxTxguwRUWUs4x6kxz6xQtfKWgkW/NC3FRFlH/XrAXg5
rHtytTE4tYptxfOfzpuw3wk3rogZDQb0FDxC4/OrJfggiZ4gFNjuFC1K7JYvwo3JZrWUu5qxhW5M
1A2qTO+5CAKuhDiFYy17rbRKpT8IiWFGv9qtjCkL0a0VB0VMtupvrdk9v0WtU8Ood5kmQqXGKBWN
1lDpquEsic7OFnAmITx60cG77fNF26b7kPtKLCCn0y97r0cX4w79/V4fsb6K0+f7+6JKqDUHF1F6
Bru3bagP0ZNMDxgeyRTOPJWor987EuiOtoGkOssHcE/IzRD0S50dQPGc5EoTlIYFdUEmziuPcx2y
K2C1QmqilaPcyBRAiJCL/gxD1cY7duVug6aRdmUQtUuDnEx4c0NDQZ+cfUtbJtmJtFUtYDibUD2S
iILDe8N6XeNtHuI1fmQls3JHXT1LC0+s0n4cORx4BmWP6db/WnyahpWzUTDeGqGo7a15p5s880Zu
jeeDoDbrB548JGeq2s/ARMuqJrOEQrZNdi76Lt5k8b/km7mL0jyE40BwNrGHRgVRbDQwROLSQN/8
z3ko9/wa3GEcG5yrmi0ulW6sPiQpzhVIVCe+WUI7z7kLd6Up2WRcqzQIamvtDBIqyFBRqvy4ymg9
lbNIYy30epJmrvS1kYTEAFgz/ES6g26klm7R1E+wUeqO+XCzMnIY8cK/2QWu8TvWr3ZkxQYwJc1i
HvZLrcjkWjFQac0Cb4yLGxLapfadg5o3QWhPrKX4OvxA8HRaty/wS5RqRBL/WNVwFfnTkBVwB5ph
CHIYa2p2KCmhtiuJONVqYQZUERj2wtZN643t7sGWlfr3+XZ3y0A+8b/P8bx7H0W0Zfb4eNSnCnJP
iSEBoFBZpaBxsmwGghs3N7dhkjeLnFRkVqdzx9Q2s+Nb6a7I6P6Cqok+FNWlQtLcMOH30+U0vXNa
zjF9z6DM0bN8LjJF4zszkXwD0tEGGsi7DXzIULxTYVA4MQ3jtRuyLOHvqT0FsZJQGDmKVtW+B7is
rtm26z/veO1lfgOKZcROPvdCj/NLqh1jSul4kRFU0tqecOdjnvzxx2wVfX0T+vcSNDP1HO2wpiYR
kxmr//Cx1eH/kf8H42OYVMgXqAxrDYIW88UCY/isQpvsZDX3DAO5gXFvHrjRJudlm2rtK62VEGOQ
uwjV+xw4B0mEgQcjuNoYaQbiZtOqhGyCbyXI1gNR0v4HZ/c/widMV4S701hCGeBmrkgrwXcE3/lr
KDNz8aXPItwkKjvbtvAp/i3T11LzeQe7pV6k4/lvCDrHKTnUNdUGyabHeLlfLbonvRa1NG7k62C0
N7bEa6ElH4d+WDm9lQQgBUYUD2QAxIyPsX1lfvoz0KwP582MkS13NIa1CWA7zSxVl24R6pepZTaE
JS2OzVPlMgcV8YWYR1GHSnhxZhW7j5Xof1Gq7X97ORqYsjXFM1qVEmjtTQKh5ifmOeRdA8yTlWEt
8tXnwzB4Hj0fwwG+QyS206TUXMVImkRNefHxrxklecKoOK+kHyzW8JoW+VQdKQOs4AKGMVo5nVMy
CqsuBv7r5eQzf8cEBU+T5z7FV8BQQ6cm9FeQqjzyl7gbcHChJkCOh8Fmg9tNulB+Jw5+c+IvBeZf
FKBbkZxPlQt+VXe7ZsVxQ1FtN075Q8YKEImZ/e5BCpcVz18NtGkoPl7apWzL245ccN0UCF1X7wO3
CSUuBkLYw0cJAujj636h5m+1bBawvYD0ILrD29L0bSyiJK4L+R22kgyTQ6Pc9WcOSbxSLAfUToe4
Fk+eDxgqzgsk8pEeQoNhPvQ6XYqatiu1hCRj/GVD4mLGOq+L1Pc3aDKCzB/WfeogtUDb3bgkSBPb
6pE+NMYy9FO2BMtIuOaDhqbsY0DtK3KRO72O6eWsKfy8AyodvUaW6v3RqNY3vgrDUIku/VvtQQrA
ZqRV+zuNFHHTOiXbqO0ntZeen5ezrkFOMnNsuF/7BZ9nLgdQ6KtIRLFOTLQOhs80Py5XMhoeAg0S
b1p8Ku4OKZwEU/8hSl6+C2X62dAjvD+s78Mr8k8pVLYwOuUONqEfNtIIVmM4W3sonzLXm7dQslk5
smaOqTnArXJRLHxGkgtwgI4Z/CJ4Iu013z0ZV7iYPaMgWuVwQN7Yid6Zj/GPhcFJJNZrbNhp1c1R
6lfsc77EnK16X4uaRjOeZOkGf/4i33ShOKJSJaMGQjs4qHSqroX1ujTxYEqniOCL1TjNKTdH2iOs
SqOa2e/nvJBxgdasHDeE3s1OWdnfrSdGK/JFBo80M6t+UiofwzjRFSm7ZPb74+73GCcU+W98ynrm
LiwEiY+bNTW1BishPnYxsoqMI34iHQrNAHJJ9Khpz2v3Oym9fRbar6qRhKJiXcbLgnR1ltQZW4N9
yUCXdxDUnKJWVbfg6F1qOGeiaeQIRsA9EIrlqjLapcWsLxKWGC689y879wtuxJd5e/LzPbpENRP0
j0SctyQgceEyll/ltbyi4xnyOSvS6O3974IynYLVQpxYozk/UcsbRCJq5nj5nb7Ljg6a8P5s8Yqs
GCuOgqs+c4U+wzQPs+6EwQqRESDoQSWibaMHGEU7M3amfHeARNvItnlP++38AOX4DcoWLmt+VCOH
0RaOtAw7B0PWFkwCPBR6TQI1CvmLdgdodxlcBADMs2od1VogTXnSC62m5kngRPMz+6HxvRsojY1R
cjA7Ga8DDYXoSzMf2h66IeFbgQMhyx/bNnww7Mo+HypZ06QhBLbb9lM8xEcXftUWc8wArKqG83wn
E3b02yaIjweHSackOAsd7WiZFjDye/ejGr/T6ltjhP6CmPWnScUbQV4syeay9Q6csAjhn5Orj36Q
2VHrAjDJeCTtuE6JOnQZ4t2A98PdkiRMSt1x9QdBpylwdr16H/HER+BVuSeIDTTCZWAuKDTAR+WA
JXSHdpIGF434oYuD08hxjy1mbMSj1N7rFbGaqvDQ3p7qdU0Y+kGsP7ZF9I2wTvUo4CtsngQuHGqK
acSArkcA768C/FK/5M7xjwH87qMEcCUZ9gwsUOtJkQ6DvcFcbZ3JM/3J1S1e73/i1G8RgvXFEdgw
SEgVt75xv+P3S3gTYIFuUedyRlk3pcDEKK+3mAiHvVdGpmbkJD33Fexd9MoWE3NQ5JRuJQqiTTwI
N7szqcMXpmkO1pxWSAQMDJUGNWfEPS/bt/EZkpn8uvRaBKUYRU84ymZLgMEXknBu9nfsmxefFfxZ
j/s7TH4Gg9fsOfcxPrp88Yg1jcskYAbYsstGnltOKdWDbRIhLqE+9Gj9Uu2eEhBz3ox9nmu6P++/
81txprSa83YU+v6kNp4rDnuUhx2eLgTeAYnrxuAwe49aRFMIU7lqIER3BZYvIbt9PaQ4goXG5RrH
GufJbrMJsdx2cmyjwfKioCCeubck0BtOd7OPu7nt1R2pSXg3ltsHhrUZMnD5WDdujrec6pWGS1r7
y8x8IF6svAq4vIfuAUb6zo+vYLjDetUcMvSAsJY4vOvAxOkOO7zCJsKRRdr5kqKTC8jacUzZI8Uh
uIqKnx1Qv4/upqPhp75ToP8ZokxTAOxL0UpohqQPeJdW606A83L2YYyqf04INUeIVlR+3J3JLzBS
yaG+bsX0rQAdnmGHCONE3TeMdg9pRp22VpIkQTEDHfTu14EXz1XqQhotzQVKUUFl9KAGP+tVc7cD
ODyhBXIsvI8AcTDWsH3z4bIro6noVikaS01arSMDH8MBwBnTp8rKpC+VvELFAtU9WqO/bcfSs7hJ
zSARM++kja4h7UYKLvpZCV5O2d+TMxrvTVHvPgyct8ZhZAXI0rAGHC2psIvNd1QB0HnddAEO/1oU
MpDVxEn5mdEDZTqCX2NMgBPf/kjcvH2+ANCgYsRG5RO+ssNZds1SxK3QhTW4pvvhbF2CAFouBpf5
QWKKstj7g3/rey1ey+ot+20ncEWPUDWOT8ieayLcRMZCriLGqNH2fV1PPZZTwF4I7XSKik9s/5+e
MmcH5LGMkG+Wz3gTpeqk32h/ewwtqdDGGSgtR3JeRBWAqXeAclmtEk1NNP/kzQAaVS8XvlNWwu4X
pk8JFI8ARj1wDUso+JT8NA8mJfo6Q0kPMbmV7pp5x3fdP1/iVJYax/IwJKdBStkN50WJ8lhX+u5a
gNhVsb622oT/lWNF9cRMF1oHDrGdA/mHUdGyk7v1A1T/HLpkL3L5pilPlW8um3AXpqFzJTn2q20/
FMo0NBln+TeT6/R3GCZ11+2RIprvv+m9M578kkgKFxLOzo6C7NTOsbQevZUTScVMQogw8J2NLHho
cwCpsWDoU6EJTQigq2TgCGZa3wec0azw8wP7dbbotUAGx9nEoPKvtnHr2czdANMIt+pM2q9y/x80
mleywUEBT89rwAk0eM0qzdVvqP1kvyJAA7BpxUxdvNgdTn8bnhGdRtxKzJrqNvFsU+LKNyo5mGxZ
mHUHX45rPbf4/XSrcbmnljnOnVz9iOqjzo0h5LiDqmvuKxWbtUS9nYFEEfxm89dhv30HNaciJeEz
YrRgthNnZR7RiHfuXmXmORnZDxg84WjeaAKhhlDvfmmD/tk4ygsSpJgu4JBrvf1aWrukPZWomYYA
vp+/Y9RqgN2iT3bDVKRWgniQJAIiRheWHOfvGqe/ek3Z6A5KS7MqsLFV8LHOCtmB9+7edn6HnVeT
rpngVLPPePgYoD25vdXnJCoBK0GeJXTWE3/1vnyQKTxu09Olv92rSOYSpwCdF7bqzWhHBS46JbLZ
O6sfr1D92yCB4aEkYttX8zYZANZgQw4+jJfckHL3V051KdU//NPE1RGFP2OqxBs4LFBAtINW+QvY
FWBAjq2lDPB2GYx8CIrixksu/QLvHRegPT1Y3vaePuqrLDWruZR/vFRMymPeSRAIQwCRP/qIrw1T
TtnartzlPVflQMxe5oZOs7T9WRfaILglh0b6Ogdis8YUW2zfqZuwXMvZKUf9g0PGhMzkJ4CJKT1r
9dhbnub1JHQqyyu4d3KrZ+TlJKtXFWze0XMIcQzUvlTEZmW/Un/0oSxvXadcTy5GL/pFm2HE2SeR
HVCiFZJMVwb3VvPeyDe/kbmx2lmTjG25UaRVYE1ATQjWuOkRJTVx0jMXj069E+5XEAtvDInc4/VN
x6A6xXqElEzHsu5SHjeqfx0rB20AjAkAYhy8zAq38EmCDPSUU6OJOQwCx6oedEviMDuxlCLPZy3L
RoWsz9Ci/FUKw263/J52kKe+ZhEERqDUzBaQQeLhsF71OHy1Ol69FIXBKiHVWG+WnPqvfrN8kt5Q
FI5aRXDhb/SlnIfqH5kTGsRY6Jjv8XAtsK0wUGJZOTwTgG+yyXfLA9NIMik9y07yuwOnJZozPyjN
R2cLjqXYfnm5r/Utsj2ZiBYdCe4C+igkym4pA7+phxt770BYaLxv7xvPiZtoBzjOfm7GN2RakWha
cysicYuYXmA6sttzEWYxTseobS6BxZw3vHQPO4gthGDCAsdErF0+zYHQhzD0OY0Xf/HxScTYdTtz
42BpmksQDMzt7JDRF0jIJld57pJPICrmFPh+giHum81e4dVo1dKjQ5U3n/PtZiyNt5VkKuAWBms3
RFxL04t/6fopWtad8KmUzG+8rjTUoeM1pBYaZyYf6iy1tSVpQc5DeCBx/a6dbgfUkooFLUL5ef4e
uX8UpX9yDotg9dnaeUyXxedoQZPqT4dZ6X0wyifirF8qpb0iy0r6NZUWSBAE2xRn1QacLsKBRGDi
iK+Hei8dYbEWlUD9AH1dKkzNNYc+7iOAlRPn2P1/pDzlSQp//7i4SUY5Oj+RSRIfNyGc/zqKben+
y0BCK2ZRfKI3CKkzwQc7HVPUNZ4fIK5HU0kUNMcY5gd7oD/ouy86OyZ2hw8FzvMTrNjX8inc8nVd
AYDr/sk9LThGYuX5hNxXxjboodsIBwlM9B5QmBPhfFOHZV1Dip6xHj7gQghwiTOUFEOdbgPSyIlf
ag5YqH4IO8+bKint04JE+jo4fom4VvlyzQKYPiP67b33j+7tTu4uAoEjnGVWBxGfFuX0wLPvKWnf
he+JcsmQ8Pd3bonZ1rMb7M57E5qChUYd5GSATTmE0+/Zwii5X7KyBZlYAgSxnCOKckMsI0B7/Wbj
tDEyxZ3KG1BMsIX1V0tsTNw+F8KQpGc7vjjAsj9kIdSeW08a/10TwKVaSstgLkxWimG67Mr+32iO
0Z5RaNR4Yw87Rthhh6b+gbeyd2+Mj4AavJH3s1aDaFLsRbfNuW+pZwgmySIKhzqHcXcq5qcb2/QO
JSbPu0s5QqJtp8V5koY6O6VbG9xW5W881+mB9NYRhadJIoesQIR09zwjkCmAv5+qRZPFwBSCHQmX
AtG1rJtpHqlet/2glWRRnrDLN0puNEElme6qYgW8ZW1rMOPVLL6kmNna7vCWHhVDLX+iDkA0Y1Pv
T46yZ3ZX/EqE6CdIeOqB1QEo+zYxxqaNlY73eEfbhW3dfPNrPjsIpmDH3WbcN8z7Gb5wPokirUVD
o0fPBpHVWIoEO+6zjEVv4ir7GJUki8vjeUw1tLym5ujjDru9EQlDuCNSv8MkQmdFg2JGJzsCN3Nl
ehUBOegZ990twPYKzOpzVbRGTzJDizxK1QMt7YrnzAyD+wWi21Pv5O2C9q7+W32axmyu7pDyvZO3
dxi/bkH9ppgmH6PNg50yup2yb6vhvXteYekkYwaUv0EJFLXu8pAyxex9LN7SxVMLWQU0XIQJ78g7
AhVm/GGX38PZmhcHbdcD/8KIF+feTp+O1ZYg+47bdBDTs9bDf0vsBcSYr+Nxw9nR+zMsUvw67Fqi
PBu9my2117tVcp3jF54esO5fwhTXhNXc1ybwr6au+j3eBHBE1+s52gAZIHktLq7bbJiJnHV2OzvH
TfqQQBzhy92Pr3QZAIuXsKiczoDtKCN9LCdXffeHM2O2k6I61X8YV5Y4l8NpHkFGxL51NRpnK2GS
8USWPsph7VzuWDU1WPsDWoVi+Dua91Ua++KUxQyQJVr4LcHRDYczzwcUwEiQwSbBdPlEhBW0riKT
8PPTa6mQx8iBu1TL/gmq70ziNciZjJl57ii/2P3UGQUbpVUEBovVVULyOD2dw7iXEjNGIWZpdo7S
dnk9w2bTAWaUuhQax3I3cp5Kbp5Lid/VhpC4Xj9xePOo4EHgPj0TQzhEJfXdeQTPo64jCqdWOj9y
r8nqiDMKWfOpPsGRlnO9wpazJaVYDchIY9BwfbhMvGdM1QmpEEi2mGLQAclsrQIQXm/cVG7SNLUj
m3AzfwtgHPmiaYgtt1ZwYxaCdxP32jtctvv7nbKF/iAuxMoOir1Slx7Ldj4MMVM+pnKXrlu/vDSh
RS3JqYuXw82HBU++/8p7S9JqVnEvXo4n8KJLAFz9TlmC5pEClXXj1QWcmLqpVJ6RV1HA1lu+j/Uc
O9vxjzVcJfo23hEKNJO3Ve9V2NLQwBqyP+zfVW4Q+UnGDdj85Mw9sSE4t2EcKXpoYKff1CR870gD
VrgOSzJoDFL17jRcz8dGREKxf0Rhj21OOiS4Ugj5ZB8YlpOO/y+2mxDWOPHvXN3m5B9o+1kPyWjF
cd39RXvatHw+ipaRUrEE9Whsj3fz/3m+ZhK6yMaqMXy6q5RzsQG0hFY7SdMxrh45Rrz+2/Kxe6wm
HwlY5lpLyIc1LGwDokubv4Umxg49ECGKMGLylrMmRApddcrl+tO0qFpOLN1m+dv0WEu3pPGxbJe1
JJSdX5SDN5iqoZOpPGSkjMCcVrU/kiL2Rg0F3kuIomFxi7dqzb+FkYW4WiKGWd4Vaj/smXOCpfBI
OpiLY6napT+zhQVHLZmjujzdCeYQgj74ijzAvqDFYxot2zRUJS6VsgLclmAAw5mKUZ+a7h/n9P80
hE5oyJRKGW2k7XlG2MVJiy8Bg2N4QAdOigr9wQ1riIupQkkRDKrzl6XqJg73bgJirmevdGpv6B/R
ZxHptaYminMBTOZzDiB+WHDGKOCCqgJZjficbOg237lBKG7B0+11pK7rspKps7TutTEjnvditdH3
G37CzRkbpvGgCmtsjkVuFJ9DcRAbtwmbmvttmZaYidheYzDYZcCQ65YZ4yXuwdCHQOLB0Z+IV5EX
z50QKB8dVG20ENd9Sl4Xl3CJgOhE2CsLLDM+XTKS3LBsu552sS81MYi1yyeyyVte0DXjAY7UIib2
kqjTSSsq0vBXqMMTHxF/ywJKn7NZaCqS30xbH8ASfLtKsCuQSNP7PXVDRhjoSHpPhEk6AYge0NDf
7AQ7mRK+vFOpUunlPcEvUYV2TVotnQS8yprgpn2AcZ6B+P2wWHbifzKDNnOgxYsvU7imUdnb24UE
rnh74BtYNme0XedK2/Worpn74Co+T47upJIr7UBwu05nFy4juYz2+MsqOaloygxgcGSQiCr94jKg
m8AlUKZp2/A/oKhOzDwUMQ99tS7qtdc+7z1d3LNukKsEY4tQVt5hEOdruuRAGmdN0D+f4NFyg9az
cJAuRlZIAbFN2A8ZGS9YDmmctT3ECMZIOiohzsq4KWZyu59uEjUh3djciNvbjeve4dL9SIJZkSPu
ScMlln3jiFLBuhghsqr1B5kKtJ2hSKTagzwD8mB/XFK9zv5C7ocBVjwwRzc+EonrTJ6lTAfkPFN6
HZqrG9oTKvA51vwq2QBS/qsjFk6t1xe+v0Q+ImrpFGDHPou5r/WZeMCPF5dBCsT/CSH9w8wCedJc
sMzQ7cfVhWzK40/sGCjsw+5+F32tiav2H4TbwzbsRkm6i+dQ9S0+xDwzrliTbWuUYc1aXRVHzR6j
ZrqwfP8nTWRD7zApwhTjN9O3/FQPgfDF8gGtU06s8adV2vUZ44H55KiJMJ67lZVJ3s7f3o+xZc1w
rQ3r81U6Fw3CPuuzN5AwzU6nXJ3d3QuoseQDJruYJJK32/8v+tioeT0+lshcbIu14mxSX2/cReA5
vl52jPEFII5vAmkIJECDrqTkt5RkSACvs4mVgmce1y7SC8q9g5yZsBuySy4ONIWfkT+Pt8mMtYGs
YTxObRhUaJFJU/lMvB/hATuYoarbsPNL70DB0UJ50sXuHzpssVCUrdoppKr04L2T0AdFPT8W08jZ
59LEkG7xp7jEzm6jl1Ytiq4s/IjEm9JfuWXWhAkZoLaCfJ1yPti5FDtNxFmbIFYfO6tV6Cwa6Rjw
2JZecIqkA9WBQn+E33nEE2Jko4sd+WZi9Gzgkda7zxsTRETj32xoSUoSgdZp+UKbuzIcOHd8fpSX
buPhSnxQwmVj1OxeLv7nbCExjaE5CmZquMBdyJJ3krwI9LsaDUONJp9AKhlECdkCucjHXV/sRcEO
a60rcIm039B2S6psKBLQvcFJxHGGePDI2V0ADipPcXmHs3HpyapKPZNWMBhEsOM/xMBa2Eid60FP
mA8VvOFgiUnqeoj4pnjvSfOhO/TnMNfc8htFy4EFXTo5oUkYmcu26Gm2uq7LLo4lH6z0eE+RjhLA
n2K+Yzd/p1xRs2Sij8+jef2lkvzq3zWNqUIYgI6xDDKAyge0NkhoJY1oQX/dgvNTwRrKhMjPbRcL
Izbv6uwqGTCb6FlrYT1aPQFng3s8GYqUzVn7DXuP72grNB0RUxKSnTYxCCJiA4QVFG8SJgaafBlN
kl2ZZbvNGEzfm+NLXaP87J2MC4fRo2sVD4HQGXRSlWljp/wzEt8rSKQVUdn46KYX7PMkI999oUu5
iekdybEo8VsLCabe0sPrsaf+oo1n+V4q/s02lINXl2JFihL2B7LgE6R9MmOrxfZO9gMvNJhZueRB
T5RpcjN5k8WkPnUBsN4cyfFxCjd9FLLV0fX0i5ZKURXXyKf/FeNGfxXsObuH1kEYUDvyfnv+EAEv
zUAe5KzRaK8r6oqf/2OIcPaUu3zp7TqM2DoAbL7xEuWD/fyxRSmuoEA0sS4aRrQXEc3bTe49miZR
w6TQfn7p3uBRxKfRYIuLdvX/BGf++evpxK17Gsgr18lFNI1m8JFTmUzzkkxPTasp841S5t5Av/Ao
8nIMSRHTowrVVgf8b2TUtpS8Sxo+Ld7f6TaGu3ggc7LQxATsjoTM+7THC4AMQ4sfVxiW0Vm/a+m9
dt9zjpYEMCqRnJ3lj3Fsl14i0XoiHhux0HQYeM5ga0sNRRdNaQ9MLvCVO7jsFFqvF48isZBRiAJi
spE88Lg8CXYTGZOxwfRspMK8KJ3WlZCNTo8mOo72QHfrNbNhAyDdC/cDK9V/CpqCvWfpCq/g5RiE
wYR+BV30dYbAUfdLlr/Sqx7wKvw0LTE6GNGpFw1nC/MxDBk/lIVW2f/gAFYp9ivaWNEYtHdbZpGd
SxrrH4upd038QxyCyQCviuDbmJ0HL1h2uFeEN8Z5BDXJjTctyWCCfZrig1maKB69qV5Y3CUouI3o
zttIVYdI5Xm+tpQfL7EMSsqFB5xutW+TTFJDsPsac2zJkCdyNDNTxfOyORBvAwRt5ojzxYDUdeMK
u1sHsuNS6L2W6nReOWh5yr379yaYzsDrNDyyFRdrPoantw+n+EhhRkOI3XS5bGaHuEEFsxOooe8z
LWOY2hjpqvHam2Yy9X5g/3uy/Rvn6F2lyCezBBYbBerLxIYY5rxqU+Ox1mMHIX6O5ci/zyaBn/DO
5hC6InvXPM2Yr6tsUAQb2HBXPZYLx6JKCzTPUaEIFhzFfKTIshl8UNSn23+03sqhaG8ncPvkiKcB
FUJc0ve2I+8R5JxLMeDsfEeZAEUKUx+dWg9g2nDplerkO6hEgUZ/BYr1lzne9qefrlTR5XTXtUXa
lko5Zgp7o85wCsFtRXQZLEZhRxpZttEBVNgEtBBgr7Yv6c5KAyaonPxBmGeFm/ve1QpriVztOHKM
2ujN59cqLPTjlNsVJ8SPAmNwBKnmJRNPHag2qjtGOERVa6o/A/vDyYjMH+7La2rup5RAJAuDTqZE
1P1f3tDQwaYZQ8KYCl8cbGokBgMKmyg6nskuDeHJk9Y22l28355eJJRnUNIx8yhoUQTqeWk/4YVq
4vK5iDPmh1kXg7Movcz7Y2E6j0FPSn1w/Y6jyVlain029BKYFjrTz/8GY4nMqtm4aFA1Ca28GOw0
FcFC9GrVaPZlkNjdVf6XimANW5ajyhAWZYqzgw9Kq3Bf28zs0sIdBiXeqB50FGl2+h+/8kP46yEO
+KdIkE7Wv0UDgnn5RwMlSqLbD2VU8C7Y3I5uauO6j3fAriQ0oSCnaXTj4VKFRPPZrejakAQLXM2l
EP/e8pVmr1lB+35moUbvv4yG/w+sEQIHh3/74nvMEonv+1N2X+mF+CJ5aqopGd7CgpKmoZZm+Fyg
m6le+fsl+LrRmVBEhPiFygvIDT5KCC0f2FgF/Hp6/6KAyDTy01YG0g8sgzvVP+umqWVYjgJGdE5q
Jve4DRXqYRD5qzTsOo2QGTlO0YiM8UWpLinXJr4K87mIeF2vOz6XJexY+HRQbq9nde2dhQk6s2bd
vJMQPe0mQ3uBu36KByWe1qZXOnd7pWTCZiTkDVA2lvBVy47Sn8YBjAwjtKeRnM1g5+uKU3E2WojZ
PldxJ3/jQFtK5RYiN/8EZObBvHTYt+P7EjTgzJBDvQ4iBNkaMfwva+nwL+TScejSEJmlkmJdkLs7
WLZU5GU1kRoAFdsfXNJrtMlLsOIweZOve8yCTB4OW0deDd4PFBYkNmCRMfikzm0W0ofXHpQGVpzb
sairNHU5mFkv741dI4oEHcHkdJPLJ8MWmV5qNuMJmQEA1k5Arsq0t2xN3J7sj9PpwnPN0UXugFox
WjHULAzefVU1WByGf/7uCwdSO/982Ad0o370iuhWKuYmG+OP7mXQxrPhv9xbDO7VcSx8AFYLVX6+
p7yWqFqpV90wFfjNiTaDePSEMI25TBvOLwdaf4Zirx1odlSzoiYz9famGn2lTaboOg3JCu5eqWgT
viTPwNxpptWbAyoH/PYxyOPDS13/wzx6x+hXV1Vm3lzFIqoeQnh5zOGW44LPL1JLXU9UsBl+tYbT
2emc/9irTdimbWCt/SxRvu+ig3gzuZce67nQdm34H8WKWA3xx1FEe1WTSHxex3et5y3RsRy1LqGn
U5rkaV+MiT+cO/gX3kAyfVwcCUd7a5b40g0Y/ZBYpe967Y/0+74UqxfLYHq89/5mpC+5wvNgA0k3
wjpnLoaN8RdBGMO7InFouv84IM23ZXTIQ2I+QY1Pi/M9qFlo/09pZfVd4zglQkoI7dwjdsPZez9V
+ScxeZ8HPhb6zv03X7CQZrKi3m/+4A3I1obCOIQMLWF39dJYlanBSIMv7YRcdixHSz82loLKAd2t
jLLzzKZSWeYEIQfk2vz38rUYqJAj6Hs2D24B3WwlZBBGuQNC/kjweGdA6q1ywGNbTL4/zdJxZ8xi
txCEQ3JoOK+Lp6YTwI1kqbWfBg+UZkhuK5gU3wWs+p9K4l/Q0jUpbaN37pKyFqZG9MRqnNe9MLFI
fjEWTSXRk+3zvGI3PL82AWZb8jjVPTw4gtLMkNIO6wnUW1VSvCIu89b65PAo2+xZmaJI8T0gbyS5
jX/Qm+K9DN23/joGYLyS+cZZyPCRhmbFNedrNCsiOHBmdwoCrwIRcKOK6JFtPR7e6lsULGuopMmy
Qsm5r458Gn1WqAooAe14ewtcn3xpW4t/Pr5q1cF7m3BRqE4YfUoR+ljIT/9IFLui2yvzm77isUi4
NMF3q95/fQ0OugAA+FcG5X76Mq/AhJiPhiMqHad9fDJqSY2Lw2Hlr7pbjVyGCtlS/tVJ0uLSI0BO
P6d4OEfqci6c6q9+Xf3p+pVRQxGZRpExaL37Elrxoe3EAZkaeHHCJtvK6UqXm2zq5ee9d/OlGO4M
H44s5pufWjAgTGtR0pARQWzomlggEe+F4yBm1IgGJ8oaAMrNi8Q7Mu1UEghPSLYsYK/36SKzr8yR
vy1FfO9+hVLm1BpfxjdRT2d5+lPLwq8n+xafU2E5u8XxB7P7sJKD650ncrYl7cAallmupw+l15Xm
eYMrhUIW7uKw1KEMU27ucNe/a4Xwdv7QZHMCeW/x2o89EH94/7nE3j25/zgfAPBl/MyjnS37TF0N
KdzlXnOfEGc+oInT9diEGNoacBRIgOtryPymvxu+QtT0eU9tuMqYm6vPTJekCqJ+6oNlqgtptQOy
DqX+zeBKiyDwURqcymcRPiEa0Ru++jXsJwB1AIeiYG1PpQFtAvr6SIsjXx4cjVsALB08xHIrsLHB
Y5ov7nNZ8+H0qbQ0cwuOceojQeRfikwdNaqtrRBqnbQMfKdEhjsefH2cuZQ3H8RH2aEEv5ZPIcV2
NloD/UqBt1r9H1yHEBXV7bUUlzT5dsvEIxg0lE4IIn2zxZI81UKZ3AoOI0qQDlO92M+qBsprcT29
yMQd0YXIA2EUkFVzrngp0CVArGnDmW+vTrE+abD0cQgJNxbqRZVBkdC5FKpWKuJUWuFbXlO6XKPj
Fg6a/Q3RW+4x0ew+/Hbqq8cEFJQ6VpHKOzliD1cI8pPDb+lczF4RiYcq0GV0Ukf+F0l+iYEdyZm+
K9g4LmLpUvSpsygUu7pKCujow3g8t0VUze009PZHjdUGG4Il1lImvDdiCUQD4b7gMcUyWH6Dw87K
tvnz5Uw04dTRWL7DsuOoAXoskVBb2fs8KSCkn9CrQo0DMiKJDs7+xN3NA7i9iZvKtRyqz4raZzqN
1QCPBRM91XlI3/oMkDadSMqWxw4P1JtS7T9BxTDzZDAqHV8bFN1sHabwFxAgalBZnikSwd6gvo/x
NlEk3PaziXDN8aIz7fBdhyISb+fV9Np21a6EPtg1/fHBYa72kEB62HU+FMqQ3Vdt7QzJptHZmJMA
lPVca65myMlLqZfvUxYLnEr50qMd7bS/Kv7OICFh1bs8r9LSuBeheujf6ayYjVAaEFfJQl2C78VD
DoF6mBJyGHycuhjsu1OKHsxMnB40bElLHWQwq/XB0/BJKYX5HQHanVs3WiDnFEliMKzUVz8PAhSy
97yS1QaFjB9ezUhhTpkZpMVgNWK04emt5fPdIpEyXZ/7lZUD7C08X6K1FbUN7wwCp27+9vgn7evC
xq2rt2e3UEaK3ydHlbr5SQjiUr55+5blOfg/k6XAQ2i2MUr4By06q+RiI/3ZPvjmAzZ7koZ6CbuX
ydYg4XkW9JYoO8SVMAdJyAuld5kqLXzZdhfH6P3Rf3VOY03RzOON7yZ6EOcwbd0JgLt3LWZoAy73
RWBxHOGhlCsjAscLLENclO+DXK3QDeTjNOIWSHeeYLAKicWkfsnwb6lUYpszTFOVMQEX+4ChYEeH
TPw1ex+Zxbmtv/HgirheXuvcL/5Oju48WDJsfU3hL5ANIBtJywbxdihgjp8/9/YHgD/GkWxYwxTi
Wn0vTTGzSjQITTRnSo0uQVXSG1gj+meoP7t9mAxwHpV9/tITQldKb5LgHDeQvCYoPO2OkgIJtwLA
sk9B6eBPpAlC6OwIy7387U0RG3EUlBH/LKGMabFKjdgYLwWjOLRe0vshytccEMXFPZs8RUnkyl3d
LVS4QBD2kTtlbdg6K8B1EBqwDNQlfSxMmIBZWEJri4OxbZ2gRIER7GF5hIff1bHYjZJSg0cQCtO5
kI+1XHPouKxe36yxprTsviOtpObcqP10cLzCN4NbDEljE6yS535iJdEP5uQERXVKvzdB8kNP7F7p
nA9CqJ9qlKE0pIOBySrGqSVpY6OJCNKurH6BjgbiygR7SPT8Dxent8waiAf848WrKE72w6VHGieV
Xib7Kw2SsoZ3YzkMT0pC8EkdVG1AQU4cT8GwRSfhR4DjEMpY9LrnyJ3w7Xnp0ZNz7FZgz+7PnYei
7vHmPvecT/ojqQ13zSPStsAV/VHtwQC0yumcsx34QoRNzVgcFYycmRU2kt1OSp9xfC6/WVytbBs0
N1WDTBLotvvU2U7JrjC1Azv4FClczrH0PP6hM6l9AGsTZRjboMVXdiEvkX2IGBe6VjNB5CR5C+Jq
713km0EbJPx5k1Mbh5If4/UZG7AY2+l88ixFgLeK9yuqjxRCN1ChoyWqrcSkvD8MRGgfmNhCTJXy
mJITTdSL9B/M8yfdSuMHJxwGEQzo5Zdl2/WWIfFc8rmLCXRDoG1xgpaMZS3eYUqkE8OpGdL+uRZn
A0nOhoouvzoCp0YPGtg/FxhjHdlMQT93x2cToYJoYEy7eo1mixwQdxfkNQu2ktndngIujijGuINV
4o1alCCC9Ohxm3ooFZEROksr+ysFzqOgjJORXZhRImuEtgxFD3+Cuja/PE2O/yh7Xy9vQfhLV/23
jVmC6ALgQGkT812QO/B0iwgO6zvyVXx/hqh7ksVdWW8WzY68hO4wxNpTLNVJ1Hg/Pae/Vr/ZvfKW
qMgGJDAgTPQIYqKHSGFWPgfrMK7myBU0rV12n2l7z17s1aGpa+ttTNyf9XAtK1X8GAd2FIqCTnWL
TMrwUIffkfU8nnx5UST4rRuSMUJQZZC41Ge63VSHtVioyB21WBXImfK40o2botDF3k3lSE5g8m3Q
d1kPOPr6DzX4K3/ZgYGk6mPLb9KHIJViHAjz2Xo4cQX9zaZGnDWhmm1H+2IuJLtvqxlscjpKxl7c
s9DF4UIRyDHmvI7W25e9RS9l89eao5CznEkpkZupDa9gqudG81H47wEaNxVkDgT5nAWXbo6GCyc6
6kTU4HpBhNg9ZvD+0TyPwluc2AS1iX7Dzj90Zcvg58oHOXXVNi0Q2m30OVx0mYwVVCi+FR69jNZk
V0Rcuu//Jnl6/xlxBzaj3O1GSrHLuj3At7orOo4XZgEnErtop52yXOS/qqQcb8diI3QJFyuC34ol
WLs92PFPBxCUL/4nBEdU/IQiHjvliwo5gckOoy58Qz57o8VVJ9zELZ43TN/M/dKW8wo4vW0YGvb+
4DlmcY82/jThNbhRmueRPsP4aW4kUOZRoKmKEqUt+TiGCrPtZ+3NyXswy68OPGxdEAC/r/85I7ig
KvghVubWT2d1TD3imK5IsSYlv2Ttw9ocgxMk5yBkNJZfbfeOrxB2vFn+IwmrQ8A03IhE0tq2mN/l
ldtV/97uYVRqLlZArUXySdEbRfbMRrBCxcVADZe6EoGw/LNDZ/QSBtr2mBxF+mhujWqXAOlMq254
HmyjtS8xKC1coRv9U8FJashzBTugVluDq4b5/caOVG5o/70aiZTUHskuUL1ZoxvN0C2LHakVQ5EV
+6FWWp07vfhF0PbQligc9g/UuOjPr8Qk/jRutSzVLjKdOtkpnJ/BHVMf7Lwv5c/zH9uYHy6ahm7U
S+01KlCHugjRVswHYMNjp1XHPgr0JWcXTpA71FP+WCTDOk/cLWeO9KWtK8nRsx8SrR5YRh8lXX8g
z/PFw2hGp8a33NpldF8MVByZVLr8753Ga/hmgz3DnIIVSz1FpU5HuVKz6ewaeKod9LOVUulrjbJC
wlFxK81w9Xmm+h4yrkf6Px6OmB9ng2Pcfeb4+SVFX2Nbg7PzvPXeIlacsCLRNCy8EdOLOVyjXj9t
Q1mXiOJ4KJCtvVD9tXEU/gK9AXHm2s/1ZGXPI3AyNdYnOV2GPgeJEP23Pec5tLhTzWgghwU5rjKj
4ifoNGG21tdzhu39l5g4IFbzbSEWvtnSDVTc+YljKBMx7eu7BjMa5cOpf8OF3rsnCtfP2d5hBPBP
dpQmU8RlmMtQAG6uhU7Tbiun2gIKWoOTwRCl2qNC+pSHS/0SFyZOZ2JY0mazQemZzjPLF8CUuuSZ
wzad84oT/CieG/ZTTT3OVYkO9p6qyd2JeMu7BnxwhvMpoNmrDxloqR3/HIskseeJ3Ampg9vKFLzb
WstEdPUrlZ4qjji24I/KYJiQAiVTLhkJLNLF4VCgVjA1GCrn/VvraO5YjjAECYKeST/eNUcLcvLD
r6fPW4kRTtl4ey+0IZiRqaf6nos8M77Vg7t9AX4vzGcBhf8FYCRhNfzfq6mLDSVyFR+t3uu2HHvA
piJ1nvWDz82WqyYMTY48jMhQ60twu86udYR4UpWX+vBfc+UKc4d84rhSV/tqKxovQMs9ecL00Flo
njlPC6rx/HpoGysdXcaVxK9xfLqx0qKHzn8NG/Ace5j7Y0y2uIUFI2TaXPq4VIMlAjUTg8QJ1jB9
ejaPAFVh+wEZdpDOAhgS5aMcoPI2HabrSwbnnw1H5OIIImWcuJbSVvaCEd8z/EsB+2jaq/x6xZba
8jRGg0frExx14bF8P6oA1qK7O2RIxV8EIwCDO00sz5FFE5QcjCOetTPXydWXICpq+1ltl8SkqZGw
zGZspYkT10RXBcpJCV/RQ7OcrcwyAJY0qlO9j1bOtIycRo7phhysHC5g4eWEO89B2vh25/b8z4BE
QcWb0w1Q+DBEYuED9814AQ+1EWh//72On+DF71W3C/Vor4y6CORAAiMwBq90fpk6g7fZStYIx60t
h6B4PV/g+VbTSRAWHYAJQxDHkaCqUcIq26GTyGpml220KQuS4rlTlVtV+GDDxKO0TU7xKgkNn2hd
RXe1zEfXpkHCkSFGbjZkEct00AAT1rk9vjuZkg/8fLBHgh9bSBlkRfb+4Z+FceVcEeenpDDwo9Uu
jx/E876e2luzZm7Rhnn/qBOwVMRJ4pvqVx5op1dxqhDcmKWrp+98vKIRux7mmU8rHmpN9OqmseEK
EggUjwCDfOQH1/FvceoM8r1j+b8A39aMdgTyHoTnVVIixxwND5dYqY55j8C93iIYcl7jCrgmKR0m
TzKswme1ShoVgJHj6jwMUDG5WAwv3p5NPBXWgCooZgzQIxmaYKWwrM47NFpLXOROcIq9At7VTzEo
oeILC25FFIWBE8zq8xrJ9C3jVg4yPJr30YN64meG/mu0rSyeziJnvg85eK4hRedfUI6aZeId/dtG
QMLFb7eBdlykBSWMv/s86PUo0mfLx3Aj/9ch1yTOZ9TFqe2cZ/pjwBav0NYI5ucRMWWyoh91DGJg
MM06WFu0y8TU5HfmtEUAyEQVd7hOuaRxhJ67H/KEGluqxTcBTO8wQSzlnOcTHjlROgqX6SxcwyYG
dD2g/BnPbtznOp8cSgu0TMuMMpHG3k25tMVlweO8+5OR99qry13dYYnK9W2z5hHzqUfkVUHV1Lw5
GGHxY/9JNMevrHUQ070vAL0yO0MjYi1+UHSRgVAZK8YFHxRzDz3hKplgrAYhvW+l+RHtBxxStvGN
wdXwNOr8wXKPuP2Fnzc8v6q6I2u0wVUykNH2US8VI339UXWzjV8lqL9x+/Mu5mgufc/dT7NMxObH
o4dG8GwzoUMkZwE1tGK6CSO/d52draV+4vBY6Tk6Gv7u1idA2zKrYYVAOzt2b8U9ZRBbODjwIE2i
gWKFJE5wHoEXhE+LlEhgdLleeGI0LHfL8p6n6L9XAkPPV2D1hXKKgT2fnc7a/fpqk8x+r7clvCuh
2ZF8Zw9r0yJwZZ96QIk0Ri4PL93ISR5EfouhpG2B7V6JrBsKB5bc6hYb6FZ00chPgJWFfj340yBm
QSLNlOCgThMnqjCPPsidMtYYjCVFyRid+qOB6y9WGXLGdaUlvxHl/s1IAr4Jih8ywnWwmy8/ILyu
iixtPpgIYgB1UR+iGRxWKLVTQDQKfuxt9BHW01qvt5fCllXKlH5QHJREg4j7pJkppcNoW1kKlO5w
PKMKM+5hRKv7/kQyyMi0UoPoZqfMsWI1ohq+F4xLpswn89RppBqPaEdkXA6k6dJhtV/tRR+gGeJ6
h0SxoJ+UQeoVIroVspED5VyheXA26mGDGi2aja0s2eIIPPN83L88C5hn0F8sCo0Kv+FAqn9MU4uw
Bdny8VpASaOMCgxg3ZI+WN+OTKDOcS8837Q+7B5PnJHN3N4IyPJikhZnFwNDkYe5zGHwZFdQe/Oh
JGmp2tfJ5tF3SC+zgTCBXFuAHV2mIcjvx7IVX2crFF2EGKJJixTeP5YruhpCupRbwIm2Mzhlo9FO
DZwvPX1Qm1ssgzbfLIN8+6GkEOtoo8iVJaMx68IO2E3RF6rltCwXeuBTJ4PGgMPAa7ArjQIzswck
DEXRcugibbmWVA6wBx8UuhGO162dIy7DQx0wUaujzAgOY35LIsnHrZZFgKlDsgkh3TOfwpFhmqov
I2y52D6/bcbp5/j8YeiDxQuAwwPKeUSsxGtqLwfPQOzwHVZ2X5mWG93WoMm7UIYn0U7+LR+wGXT8
726AVcRNU6PalRl/HlBghh6YYt+dsPc2gd9N78Z3f6P+B2XWKwGErG1fhJM4BCQKrYXsHrp0Cwze
8TXI0ROyhDAWrdTKY4QEP9uMc3fz7tzdJbvyxE9rM8vT/uHeY4AE7Y7X33IzPtXM1e/p0JtgwBFc
vpDT4w4Qpb4MvcFNMVFzU8zsooiFB2RokhPyK3s1pYj3CvFxtF4iL9zrrku9senAfhDO5MG9qEU7
aUjuGavi8XZcwISLHKtS3tcO8duYbMKbdPdd+GfJ/mpTUXbkqwsMIRdCjk9ec0z7nFB2F1Az466d
WoBfQW15fc+x6pNQZlGSVOvFkgKEBrwJoS+/yQtCcTCBVqvdiAqTyUr+7BjW5YSAVfHix4ukfa20
R3vMhA4UwZUitKWCB8SsWO2yBAY6D1JxckGDu5XKQKav80IkjlLyzYaRMqULvOOz9V1TZOGykNpr
6iE6gzG1ALdjMqyd8Ujjq7qulsDvmAfAREekZqI0FqH2U2u6SysTuG5fI9R+IKayfkXEKk+5kljg
gRUrEzIfa691OzcW8XhhcmMZa8sayGbKqW0hAvJC7MaJHztwPU/clQ9xX9Cn0cPv7mo2g735nYO4
g/gPJ+dYePBzPr2NOwTUtHv5bCdSsRoemQ5tnYTIHIJlc1bjAIH1F7NelM4Fdkj4RVPNOnLT28kR
Cu+DKYUaScNdpUXdYv+nWUl/n0IJguTXo/KoC+qul22jPIvIil9WtxcdhL+m9TuTP7Gzl4/YxAE4
3ocNDs9b+HS0lVDjC+EgthFjaRSSfpiN2BlBIPlmsgmQ1eo9flkPDZBlJDUe330q6nIPw4I6i92x
81CGat0GQ/SN3XQDJceeEYuuYrM963Av1uuRfagoUKfAlNuWXl5myAu1vuOGanYtQDKwk4UEy9oA
2OfOnxtxAodz7FgbW+tocr4IztbLcRcMwCeRbMyHE410PAYre517zRfFCL0TKCj/47bj4Isem+xs
3T8N9FC/iB4O3J9yjx5O6dOPhR8ZGgiLtY2dpceRRLkKeBnoiyawLoWZsz3tvGC9Vvo3VxNGGQHb
KxjI5rT/Te7dI3u2YT7zazoqKXENYqVL+fqxv2VMgbKVPdnO+BOXcFBpI5uitrZOABrA3JlQc3wS
QLEhsOg+RrV+u9+y/thsSnlgr5u/ppjGmSZluUeVEhY1tL7yETvBOyGgIXKkSxAqHT1eDoSkfvrh
CZDQ9QugWOIaH9Ub39m1a9/bEUEkPaTeUJdtd9fZ4QiGfjxzaN5Q8KDrLCgBCS2F1KFYy/6Y9EeR
uAnnJ7YmbnlBY4n/n4yRswY/zzlBLdPHHFWxgU91cDWIqUKUwWuRAL/Mcx0xRnjtcW9cDUMUMPo5
go3yO2H2I+fh19nvqMxLOj1CsxCjM+DEc47j48xfyPR4rBqarKK1i9offP+PIdR8SZ1a6vNps+5n
K4GvitW75bXSopJTdfZWCji/EPpPGQZcqvrxtkGtF76dFq+CGguJfD4siGE+oGba+KWkAZE82FhG
VHpPKIvfPLmkYttAJEvgc0UAYI1Axz9/JchCbxfOC5YTlxqgnp/LOZn010z57JwLhBgDyZY/d2+3
c4nEOCetUYmjC1K+QAgkUP15FOh/C5LGFZ+Q8U8IStKPFsyDe3FR8ohHsjXmVY6EAqfSQxZpgvSL
tXMtpJP4oJDinLCwMPIyattO0sqtxhXMO0Sh5ReAgfBq7w3FcP/hSzFeHF7FFwvfXkawuACHpHgh
nF0OyMx3xH0NhlD+djW/gyL4Zlbmpq9paqr/yhVlX/zWiiFU5mr68wPCfvnbgNxiYHwoltQNmrSP
IuSLfiTsLDZ2fXvMv+M8KSKo7qbjEx9HOtUgSoTxs6ebNPmElYMDIGl9oFKm7nqRtHuz/NU09Kj5
NaqQjEp53ZPHF3tpw1M9dDJwe6OBABEex4RbdDyTBNuZ20YlRHoNw0+Up2RsDyjIbpByiBd3prSG
fS3QL4IdtYK1+7Zf6XcUa2NnfDafjqRMKDORRyTTauuiR/ShXCgTnjU5/uDATU/sktQex7WgxtQQ
YmfbMKsVUQc6VqhOqvSn+DUPJMPRoiG/+IBJpnfr12CalStuF4ogh5qneX4NULUH7xFju9DwuG0d
erSX2p3UEGMjdeH6DDFsjNTvSt62KFnsY1jGgzo5EQB4xY26VZfLLJuuUZpXNQ5BDvLOpiCGxFPu
9HP10CqaMjVCdC1SmfV3JVDdfmDRxj6mWiSJDc0ta+SPPuPH5dsRvC4A/rx5T4AvvqnB68i+1Hmn
cfz7LwIfbd2E+3Eaw6/kmv4L8k4rWf5/5R/pd5IH9hd8heJNQZM2F414eMCrvzZTp9lhvpStp9nN
u4+ZzduM8CGXtR62kQ6ReLpafZ94otLgQIjoQZ3pb6lJaR5E/CimZzZ8KP3w59cF6q6uLEdGZrZ4
9gIY5UDWh0+TYp/DCzpXKfP5VclhXHaJx2GLGGXCo/dghu29JKNXP+//o+H0TAd5SwxQhlfWoF2m
qSGINpn9Gfs6B5cTM7VIToJwl6bDXM08DeEq1UJmorV4Y1P2WzJSMu8+yyU9lCksqkUegKQT0xtf
+y/nsjiYCRlhLX9l+YLsAa+axhgyM6gEDjowPwyHaKduwL1h8kgjklm6MFCEAyEBIp+P9+hMgfmE
B7KM9S214D72MzlcbogmwE9+CmPlM2rPEQx/0V3wcEgYXRK90vZsVySBzbclWY0XYm3UIEC8RI8B
6S3L+Prlv6ZveEntFamTAz2gMsK7agrMCkd/ncbWSeYMHstiXwsN1J6hnAjDhfKVCChqFc5a/lhT
15hUI+GMewWCfWb4ZfbKI/qfuEynXo+q8UqEo+BMhphZjqGn2GkGd4PDasxDM/tHy7usOXyI2HJW
AMTnxAWrmPlPq7e+pFDGHdfGYdPcSOstwDN7Xm6U4Kk8VpsBL/B+p7KG5TOuQhhZbv0ali1GmHhB
QcMWD5yZJ8PgX4+f8yFd7tricLR8AuTBy798uFKYq5KUkKwg+TalwlSolqNk16ROywnX3VaOFKNg
a1VLQzsazd/XJHqu/oNZYt1WEkItQjVGhIQZu6i7Fdk0KQ6mjUpKCwBg5YtqMv35C526rEt/Kwkf
q1rkzKCOoYU48W19iQypcz7NceG6wVlj2Qg5USWmUjkpCuhlbu2T5Xq3vq0PkvIfDvGBn4ilAvoV
U6dz/bHZ9D5ntE0CpYmtVi1UZlugE+eK0xKF4C4FcgKAm7TJascHRNN0mxsox5WHdH9KxvY+y9CU
JCLxPqFk36cnKszX4NvTZA0WtJ7Z3ewRsP/mfRVqbYNMWWhAvIh8FSdAEX4QfKBFJ3/hHDJLyc36
Hq/iuia+JnqxSaDbr2VbaDYWXkSyMRBMKoye90VNJ0SNkql5nVsy6VTmCpqw+sPyBcKpdiAJzsIg
Dpo4T+pvd2Kx06B8Xro5XCTrTv+9gAeXfi4BrP3oNidhlWwzBcCxipez4lhcdbCHMYwzg2G2jyv1
j9urazMG9Yv6qilKROnHndFU9X+5nkUNGLowfjcLUX2aNWvODudC3oJiGVMluM+WOwJ8ttAyI/8E
Kwtw3H81bquI10SLGhEnSUuSZk/S4vAJ+MYsADSSwTzYtGL0Mug1OX9215+/cf8cYdKGtQyeAH65
thgkmMQ7g7/xnIgfEDCOaaqEv/DJVFLHgKmWuP71mfC9NWykvlM5S1VN+pWQjg2VJN7bZt2I9EJY
gF807FcDlLC3Npik32ujVwXHiPbQKuoqHE5WmccO2JHZ1Q4HQUmDjM3ucMHGsDvKy9WBoqnu/8+i
uN3oKNObvD064J+iq6Qn3Vv4q7ayUY00f/bDE9zFzdPAFQOciAtD3pZMP9lZSq1MOGMhszsWjjf7
eTBkfAGfikX5WcXB/O4CdXPOkYQ9h2j81Fc9jc+SIDdCf9i2ZS0LnJ99rnc3o8Gq2fs3BbpQlV2z
KJPVVkCbVyUyDwvwDoXcAmzNuI8JutQaoGNhfIkFZSR+cy6jo21OuzOX3Y0g4IwxO3HbSyNM3jke
ThYkjmq/UBGJHkw8MBNsWmMNvyZM7pLYrdjw95kEQ5gFNy1lum7yl/Jwf/XO0G5g8RdrSV6DMc6b
H4LRozIeGYfL/mjeTq25tLJiTYjZxe0T5XmgdGxVFHQmnt23ZBV956FBd8gbikN4I58AvwW6sgzq
5cngb3s9+AXgA3LAtdPGT/IZ1/sCPtrB8qinF8IJ2HOpw8uowT1Gt04Ecw0qxxSSmbctOaVmEY0N
f8UUSU3sm57aHeOzSq3NokN1qCDKSxJlg3pxX7FKYTxoyFGH2Bra/IapC/fjkD/m6o242mHXASiP
b7Y8EF8iX3CKwcDmwCWX1rv4Bjt+83rsMNDeGs+rGXHzan5LwjumNuhYX6abyVqdmtaRPMx0mRjd
H8oiqT/TflK1D8rQzej8uhlgn+V4307xH+8BkfAG9JC7hZGM4txu7lqJxqOGcZI6Mn8PjBAnooTs
Oru1CNYsvEGuynOK0bZbVrAIFKEca4e+a8DEXEf7GpbMHN3Y7bQ8cXA/YWnsMsRzqwiEzDDK4oiP
CZSbTwwk/wMEKiBLHmQE3I2uC40mUdHpbUGPn24oBv60vJ7SYdnSiHHHI0Z+1Bc9S+3e6Zrar4gf
17SYg1s4c5or97zcXY2i29L2fAhtrgbayleUehG4s+Flsn6n6g/6QITiHeLwaJJZeOEPwfc+Bdsu
o4YmVny0/CJiRJp09TE1VwV4uiQrvYt8Qh5/m6kDFtRo6nKUiBmmWehl9R1nkwgAHCj/HBW/m9Ry
8uMOEKWJpXkTJdoZIgARMJ5TIw+Eff+4LVEBPz+oCkKcyJh7xxW1jjNChrGbQddoJs93prvAZA8o
1CBxRL42mjFSp8K9C3Ut9hecAxu+NpbX5raCt+QGJZFgbbireOe8Y8kKh2LtSuEXVL9v2Mq+wiA5
Q1pbcPC9iCzFo7yEokdLiGr1kH1AprV+qf2AZ3+w+Jn2GwRzUMQN2w3LvRmXRujYsgvs7l+5iFJO
YMMm2yRjIEqfwueBemSt3Q6wKwnB2GMsoQ/YCBWCdV/pjcJRK8+5eXJpHfAqc3t2wOou0rf+gYqx
UL1HXZTqlSnQdmdobFxXTx2xPPw/940OM26dC93NaijCbY6ZPf4tA573WR/aHt8sJuu6KWEomJ85
jqtnFp56Tmsoxl/Cf14FWwpAUQyZKbPAyPnraf5GEFsEkzOg0gwfKcopM7/pUgfCF0G4mL5ZxyXS
6WPzHjyaz5Cfs3RnaQIscYK0yd/x/KLmxjFjDrFUKNNqYBAgdqZ584BGIVTdIgry5N4q24KmHSoF
Mk94ZTA5bHm5ieZSd3XiIKUSWVkorI/m6+siyGMAb7cV8ZCARJ4GMS/N2LyC5HlQwyDsJs6L4U2o
I/Y9lwlzd0n9slpJCVnZQnzcHsX12bU7sSwdu/17Q/AneOjLyupQG4h1icuxTp/Q30ChQRHIMKko
e5XbKqbBWejwvvY/6H72cVQZ22i7H5ZAlcn9VarDgufW71uNG3fJA31Iz1e4OH16SGiVtTZvH4xN
l+DlenZ4ZPTpaHScOOcujJ6chhejtmj8k42Nc6MLIRHn3f+HOCZa/xa6L0xSOWzCQWoBkte4SIHe
+6irCcSvBaeJ968scG+M1cIlU6ZkmJfcEYU+GjJRoJAmjgyWnZMv9dMBVyArakYjUGP2JlCMIrgQ
orNffD7Msd1e2FmwIzOum8h0ceIBRSbKGYfFuZqso6mxD+gXrXMKYCX2JW8e53SK4P2qVl+oF2P0
41lW7W4VB1IjcpBr7f/cax/wPHflWdSI5Y4FHpZ5hIIoi0DDLh+Zg1U7LnVJGgo7YrSyF7McPCO7
bZDcDCs/vgNRbYQxk14vdYf1E+VzeLcHLhtIp4K58vF1gJkeETmoo1wRj43X4C0NE97uN3IesmPV
8jUwkJ4zIbNpnfg9FS9VaXClgX5wKpitG75Nroi8aFDv6Euw87C6IaAEH+KE52IstHN1bBurQK29
nnR924mo2P7fOoGsy66RLM9nv3ZWy0vUbR0/O3T438rJVkF36UHUTuU8VL+6JPCb7hZrRhqkX4ij
hH1UDvRKId0caV16Cv3SZpEUseUaQSQbJH++HkHnafeFVUb651f/WbtHz3N2WM8aXIVXHHL22BuW
SZJr9NMFt8ARK7K/ZsXE02d+pAelBnq0RFrtxnkG7CrX/0OEh/2VPntkcsFiKQ1r/ZymFxXErOiy
8+3jBU0cNY/VApVVj5i6ULxcOE2VbUjsJMnKxVufSlFTr1g/DCI/r0O6YgKtM+4+JCvPzWzUKh5I
f9xtT+yILJBlyS/ReJJGcq5t8MVaQUksqo+eIrKaJwbjO66FoRSsqntIiMtLvBzWm0T3mk7qKAU7
guf37vDWAGn9GTIZ+SaqS+7w6tcvdHPZUVdsNQWZq63qIkMFlMNQb60/4ZE47eyVOWYOQP0GBHVE
GctTL9Z/BXApH/hMM3d7bYCcwci/B5bd/bMHpqC+NZ0zc8MP+eO/ULstIAF+TJyn4y8plkh3+EP6
jQnoEPznEgWdR6K/VLtRYpP2lhXCXVU3KlciThrOnHpUUWCuuViq/FQdoO2fIitTzrHKBhzZsywr
RmE8zxd18s9kKNxUZBpt77/L3iOylIGN3rJ6e9zz+/BGQFUku60uFBVQEubOz/nvOTvZbCw+mUiF
fv5V2DgMgua3/C2dUXVew5Stjco39slLwOiwMnaa6G/ae7qri/362yyWBkxr429ZgHDDiFG/oiib
OiBk932AsPWEM3iRN9dBdz8OVoahWA4FC6kFyOQ792zlFJYIkQCAHsQeVW8YgwnCwiGtTUJJY1v3
8Br060noxw8LsVMlw5G5iFOJ8c6fIMlWe3sOaKDDQ1bGC0nyUEolmrn2ABOxqSBPExhBmL3PNVMm
ZuzTCJyIQUDOSSSDitceGOj59zCs4l+3MHGte+or/ajcqsM3Zt6oEj+auOUBGerC7M5F5ELLtBvX
F7BfLB7tMyiy+PW/tnGkueRo3jCPVXmdDSt4hn9iLcnpgPpr5sAYA/JgevcSifaC6qmqAofnKGCe
zwR77kUSs8/MDZFYkGnGjhEZrnKkBBB5S1ppnZ54C4R1fGQdh74gazDZ1IZjsYE0bC5JHIoTqVsN
B6stXe4SsfiS+CP0EBDR22c35hHUUsP3AncLfmxB96oD4Oh2lGJ+hWU9c4yOqCIj/FE1h3+NJJt5
dL3NbvnH3r1shG4QVDSJhKpRwekfGEXbZLtneWjxFiWESyRfhfqVbsxlCD3CjiTN4uIWAtKcpG9I
BLbnIuKJgNRB7pIrY8SWdFDutMQ6qWm0SL/vo1MjWbujHDRSIg/aviTSFOwtuLsWo+drtP80UR96
t8hexNG+Rpxk3r99JP2MqFTzNqY0+AjYNuUPJ1rIXmijXKENpWGX6llHPycv2YCdKJgWoGZac42C
+LOr/u+39QF1qo1+e3juQw8E5YEXOLvH2+3dS6ScYGRfHmBUBCAcMbf/dwaYxi5fJhImbfy1LTMl
mYyUx93LdU4Txah9A4Ylua4J+5u2K9Xltqqx7LOM87DeQwFCzlvPRpHWWyLIlQgFvWSe7vOUq7xh
FnFNbH/tjwO0JW3MF+DrGYhfDMPhhRu31Jp/AaRK12tr9I6Vy/hZmjYSXFTCf9z3UhlUr006zbmC
nGwxoboZofMp/n6yhgBXI1HSFWD2uzhVrINKluR9IaLFGl/ysAzR8L3nfaIbRazsVTbEu1+YyLgs
jZn2HAGYbCKLNWM387mq+3EVeBK1gOCP+v4s5/rZ4DWXhPkbTKc52wg36HYRA8lHQEVFoiJLddJX
QJaTV9gvwkShS30caIX34kNbS4R9n31qCWxWu5Zbw21kIbUAVbR3r/d0xpIPkMzu4fcAzuOdGlMp
h5VL3gE9EpzvXMGaYvNZQz9MPTTNwYjK1+CWCBSnSHtEoiAPxlwpnUk2a6lgCxT1uSNoNBRUlPcP
HrZ05WgfjkUghl0N7Lxyz9PrR/AFjuAvNFN8qz2SSp0F0n5l9SeXPf08rmMM5uJ0yoN2j2vv2A+s
5rsO+z+jFOh/Nb3gblUdFbG63f7Yvym67Kdchrzy2G/wp2amOMxz1YkG4YC1vIdNxjmf1n7eFszu
mk4+iKAo4asMV8X5j+5eE4pX/3i9kj+alyDEaikgnqYPFjZ7YNRWJ0sqnDa7lrDZUZdC+l+fk2or
e+KrT0zGB6DPm7cqpg7YvQvbfZkKEaMkTFNqBsFYqDTGYnNXbokgkAvDZV7/Q6R9dHl0TZI4PmgX
rT0NqMH2KMsadLV0tzWzyWvSHiYD4iHTJpPusiZyfFqWP4IwGday3Q2uwVQVvpk8ECtq99E+16+w
acNWH3jz6pxa4v39795WMSOdTum8GKh/N85RitXhc6BrvDdJ/OR5QtD/SB1bBQTtI0nRDMBKL3/5
7PvxYK4EDYFkzfuPuBhzb4btE7uh5cQutrtDVuevKVEiOfyEpP46F/H6s0Wlt1ngHSJv6oaPsBkI
giZUEpmm4La76o8n/P/TvY4GVYpOCz6jk+qcV4WdP9sDawZb+FvaXPRgUg1MZwrxamlxOsxUbkZD
Qfb5yqAqiXoPskrpwpAGwse2LtNNjdTSsMqHCJQBo1r6TAWQXyI8r+0sTLgGjjJ3+tqx9xBq0kO6
Fll6zFHZCLSsJXq6TQPjiylifP3Ll7zioImQrW/XHEnWUICT63wXHi5sZk7ZmOVv4F6op7hX50MD
TNmbGkSKhRNLgsZxOKLadJSMQiOrxyOPtliZ7nrAeTqUyrDqGVPNdDKZRVju0EpehK747tkaNVow
p1IKj/M0Bcc8eENCuJz1c/L0xD9WlpYx7ibvThB+VpeDPLnM/Gt10WffUBSAt9i7ZVgEmwLJZuXb
ZrxL7q0pzLXwy6CwGK/A21Vx0dXpaM5N8njK6gVVhUK4b7UONjsGhtWNXZVf7AMk0WsmSz4mdRIO
AjJu3Ysf8GMF2hQsTEey8N2PsXwX1g7uI6mcKB45Y+oexMziBqsRDaMyXEs4xOf5f/rNtb78UQ5U
0zkRTwsC7N03PqepHMs85PMtErnKarPPhLeCXZk01Ydc+mCUk1D9mPAeYa0P1PSdJX2I5cYDnEBK
NpBe6X23OFpNgGFgNriGeR3A6h0EP0+bzyGwK3XHEAUM+nc+HEeUBasQ3wmtCY+XlqdHNBohoPwv
bN3XgITa5Q5PiUsFRwM89Gyhicn9/7GqZfq1Re5LdYmiIfT0QvmBNwsl679mZNlVuQ8PS/kBAhJQ
03NNlaNeCoxp1G7p7qTDk/wcOIcadfBMxeLwZvDJdr00Cr6+GZT28wFkvnOCoOgEPvDmO4LcwCG2
nfkfrPHxClG+rPUjuAAxgVM9xqBNO49eDMN7VPopSyeWLgmu04ncdx3VErWZ67FHWR6nbJlWrRZa
9Q6dGgUAp6QjU9LZkVhdp4j/V3YhYwCGmBiahxDbk4vVUP8AU3dVITnuPC/8j3NDtZKlDTNg6jbG
OMaMFK+PaTeuUKjulgcT28TtSQcipA8abVdLvZKCWyWCV0vOLL0Fg+k3Ts9oOsXDqE2miyYb16lB
P1lU+7NDWuf8w83+w4GXW4L+1baEmxWE2Q1c4KGjGLwIoA+tuZVXIKoH3PEz/vigdFXaHcplElJI
Iyax++DDG994bDtyXeEty8bDrxyC9Qn9jNHJZXMoOAsia9VwXsQpY2UkSuQBUa1dh+sB9Fmbnevp
5kFM3qOfuVNwCReCwJABW5+MxkD/B1OOH3GBkdFN84G4YBHemZe2X3aLj+j4B2e/bO92gg9lza+v
zLz5UxK8ZYc2UnXKTaq1gmgKoyf1mQezeH6EE+BarRKS36puTp8J1NAWdkanQxT6c/X6eZWFM/In
TXsHOnqRGKpnkT9PljPjCIUYqskqkL5r4O0t3/TpKca/XrJFXYZz6Y3s7kfg+PtCz6um4Ec+CIUO
X0a9D3OC01sYrIXvCA/J7POf0B34Od/C048JRqV/fmCeVoZUa0RPKmxSkZYyfd6foRXICcvkfaVR
Ss3G1ANmr0ArGBEMmIcrl0VHmja782WguGfP9jlcFClz17CbpnBd7fPeYwOVqwJNw+Fg1Qp6mVuZ
SeMftGOTtwTt1EONXt4IhT3UwgZVS1C3bFQstXJd0tV3l2KANRXLVW2oz//qaaTbxDsyvRtPeyrD
kRFM6xUYYxKUZ/ALSaDkmyfa1Q6xajKxJjxxOOaTzSg+M+ddIw1LZXFqGBVhD17reFzaJfpZ5Sv5
7l+l7DmGpqf3t5jpuvVu6+YUr2Yxo2MTCd/XxgjLoFIukot1ihW3QxLFurl5kq5F9If31wtSSdXr
P8VrFmbLBtMbWSAI8ZlT37QwP6xQuziTlEal/b322AbADUTXPwAVOTnLartQXfieTCA6rvfVBcSL
NtJDu/14yIPQxYhSONqGG1vVZGeCC09nBJdhJByghRTExy1bmk6MC+yQYoIvK+0E6roZI+pNKZRX
km5cxExW2dmtog1DiG+CJGCX3L8JhyD8MMorBPZs9Kk5u59iqz4xdNbKkS9f6mqsIgbBSF5IBY51
tciSnT5d76a9AlVuIafWJhwC/UJcH/zEAyGXwlAL7S6WtqJH3WTXHDIp8ErsU+wb8gmruWfWwVf8
pSbGRoa/+mRQWqMlp75eF0mZlx9ubEfSGw4Xb0GHBaCFQcqBypX19A7F0lz4pmFLZkiRhMGT8XvY
9S5taPSnP/jL7EV2XMFrWi4Qa/tl+uIX80WKVTBAmworq/2A+rR0pBk9BfvUCV0CjvdwsO7cmsrc
/cv+IT+JLcF32ic7aqGlpDZns2+hO1oNYLZTSyDiCxrMic23NCxqIkfV26n4W6FbQq8vIbJN39uz
PBnL2dnY9sE3KGRvde3dwa+xG7hYjeEyCrb65/cypN47asj0cisG6eQpE4b8xni7o1Wk2z0zUIcx
IMBu02v12d3EhvrKjBb5pSejzYk7YY9Jw+oCX0DxtR8Hn7FuurQ7z9PD59a6s9l0mqicRRg112XX
NgKoA7WYmd5uKEK030x4HBhQjmqynEmOr5/vFJnjLU4cm6O5us4nyPYn95tKOhqAuZyAUzyOyem/
FYXBludZnUp2/u29fCJYo55HiMzNYAQG/BSor4+c8YyUJ+iyWAy8wmxkrzFYngEjIivJBuTe7j7H
tFRKAvBUBs3usB+QcgZX/s68nZP0YG10kKN4/Js6sJ7C8N0cG9eqbR74KL4drYeCBvDd2QjMaTwJ
iZ5llLw+Ha7LvBQrZaDfUV1eLQJhGVQEcU71h6kCNmwAnwFm3QEUODnLV8aLsoiterma584Mm/ib
CCEwlDH1SHiUuJ/Rdo/n5xlaJGY4yXL6FzxyoYjzBR7lXTZjKOZtgNSWnXC9xOBAKZ3YfffetOb+
1yANjmb9mkFyxXyfeMTz4FYbdZ2VVIrKBvLZ86yHnADvMZvfUU7Ae/HANmTqLfjoiVT5KwtgmhAB
ETmxd42RxWwXKmniE++3bxHVyBcOnJsDsEZG7CdROfRQeTJ5lQfx4QzCiEaboJHdieCTIa5bpgpQ
NPq6G/B+XWphhSZCkG3MdeIcaOdeO3+d7wbHOJ1KVB6Exz1Yf9o9sTH6/UOILrscsEiyHRjS3ihH
iongGDQzOs68eUEw//OG/kE4Q0bNmE52idI7sIk4QYc9KkOe99OpKUKe3otIDX8SnvIUjGoGABIs
wknB+WfZsfNUtngCCeL1O1x5VSSw0jVWX3zKJuu5e7RrSs/aZtNhKQA6MLnyrgWb09X02W7+hVjX
FZBhIU0/STQUW2/nu2h3NMXVOCDgmC9fWfhtf1CN5oknoJfeCFvvFkGPqJrYex71mVD+KIcMzEzH
rmUNzQFO6ZvQkQCmrioBuKafrBLLSM9o5gwcTCFayABurWcqSeXftjDfI9TdVn6EyOP3NKsFE0yy
Czr0GLUWdUanFPpnwu/MBNlPesziuN56dLtIHtaDleK7vpNT/tHdVDWy1MO2v8rmE1M+h30C7Ng+
9wbKRG+K+9bu4tAlncHIL/Bd7dRVBKQyv/Qign5CFQW+66wycI7tbsjt5OpzrbToYEnzp8QkWnZs
3RNDe+7swQAVy0eUxuQMFPASAQpzhw2C5VFI4XPf/iN6gP5Kc0v2dsKVwpI3eL3xh/99l0hjIhCv
BfBAWJ304DWjoFByafBDcEa66ksSdlzMcmaFYxp4RrLonunRUJm4ZAqcRFPmofPQe6V/cP6Oq5e8
FjdNUuUa8fKLQR8/kmJJmNH1b+Vkn8KaN4Yc8zZrswL0F2PB8LDpVFqdoyjN2MyQ5f3CeaoMeGZH
FqDDBTehIHGD7B9zDzFktKKFZbT0LpLoF6IhwVizft8ZHXbuefleCkqbzl5vo3d5kweoCHgpn+Qu
X6HeO1KkEL+UB2z8DRr0yjqA5q8YPz5eZ0XNI6sJ9VX905mUVfAAXRgrF8/2o8DlYjHFBQibGJFJ
fZUxEsZo66Bo7sjdLfkjs6copE8Kew4QjS2OAhAOiMPfTNlgPpTutAaPsmRTbZp9hIsZ2ENmmsf/
Q/znd1UgbThBuX35E9W61TaaqEZXSixvFaUnRDSdyKgOUQCUW+jfR2u43AKbDKLFQHn99T5/dilT
sssZEWvYiHKrKtkGPvHUtV+KFo/lZCHz/MZUieqaOqMUboLQKsCJA43GcCV8ohjU30P3stRpr5ZR
UdWvlpynZrpnlxozugvJXSlNe90s36+zf5VdqEOYMsaEJHlTOyVlnw1kGDEb1uDuy1lFUJKROJhb
d2nUibTi/0aH1ZoFlVdf/yDUABfATLhmr546rs00A5JruycqN0opusNJYc1ZCvU/8EBd6HZ2721Z
sjHQhgTt+zDavqDv0KeFR2sAubDThWvCLk7iUQ3+9rECLVLWCfkznFz0cqow5J/nvfnD4AnHmr8t
5UskB48GbsajXWWWSds2nzeMyHk3di/jZk12eK/SGQQjShBfdlDcu5GTo9ll2qJK4qod2TbhGr2o
kJRwbCzxdnMTbxm3SsJ0FAxwfPV9ZNH8nWhIx4UGuhK8fBw1oM3HskKTYhd97OTW85s1/mu2jrI9
UyuDuaceuWrpZgZLj9pchgsovlfbD7/DrCa+d07GhZkEOaS3+1repfMHpeU0D7c0q/z1GUdJyQT2
TuggkvQXlaGZ4wgza0ZJ1sALb/IZETOt04asCzogZ4574gicI+Qz4xCsBj5xZNiK2xTyIn7P9Avy
66T20ccJtadNrMsc+QxpxpXP5H43c9XSGcC1zioLSGU/Wdf+XG311knDUznZioGH9fiiHfvoKINZ
1RNKTX2Ip3EMq3qmKNPr9HQ0xDV8K9/Irx0dvbRsSycBJwKv5Cgt3aNImi0+lloExUlG2o9y84IP
x2sD791ARDXzDjajzs+m1qVBK1CO3c36W9gLLOD64a9F+Ky4iawvcuPCvnjj09bJMrh+HS186hXQ
UzP8I2B7hfga72gzxbbtPMXooTaGZO/wb+2sAiZPDQnAFrN7rOcppb+F40ab/4aI6zwy1f0Aa7Tq
dUVD3M05IKI0mJ75Dxc5CIfe3Ebl0HorH+iacnb9IZ7dIqVK47X35CIvkU9MirISLPHrcryL6H5M
yqPJqsqLBaiNuD3OYevZVy6d2BZNGY7IePggCu2X1sBnEWiJpdakkAw27LjNjJKmNT7aND6qdXJX
LGe98yN2RuhfiKJ93dbBBQ6pNMGnFSBS3rxmztgw1/RZ7IwgFu/fQzJfrHAus9QIMztUBIE5uOD3
uul53AhDbxNTiaTHHVSE9zyloxosT/fno9mkAmNVqMjtOk7wa31sr48IZ2l8YORpUX7KmlAaOEK4
P9Bgdl2Z2r6gNsU82RpN0Z5jSgYONcO9kFYPwzVF9c6RBW8BOX5nmKyXWc0TLgDDgYmJPhzL1sLk
Ncuc+w+KzgmApKnlP6ZlSdriegj25gF5jc6roQ6J2DGHJaqroz+Ob3S/hpbF5XwzyNIiqblc+LOi
xsci8UKaz6c3oNVsBnmntKiRGC99IRPjvY6EctEFE/OIzExZYiqlT1XRyTO7fCgpaOA2V9ua67aj
FvNE9Pt7oHE+tTVjU44Dj8oNVc6yvwP+GAplHpYIVI+TfjcPhrymW70cEUXnW8tDn0xO32fD2Qjz
or4D/fiwKVTwBor+G4n+uYmo9IcxE8a/znWh2x5AQTMvjWJTi97p2hbDkMzt4zAbcmJTWYs7K4k7
L12YG3dyqrl1hT9xVgkkVgrjsUiUofVe/Dz3LidNcVwU0PwE8gYPcWBRwWxDXipTLu/YJKhe2sre
BXjJmJfEMnBoq18K0LTG2kQwYnXU4Mr1vWY9VQm9hnGHn5O5MhVDjN0a5vUJO78kbSy4cLa/jaSK
CtRUOyefur3hfPcVTkS3OORkZ2kADucHejVnYHtzs6nhiSiwwwzgKtQ/UBNcJBy+N5aNHuoAwhml
KEbD2Xo1EVYGLWGTtE0MTWaPoQUll8eiBoytw8aPdhJ83CdK6jbAcdxgplpYbfMfimUQKr9VXvy7
I650ITkyZ1tZYht+wdB6y3srlCAAqDBBSGIpnU+0WQ6J+ANS53euI/BNEU+nMqjuUyRHq1LMaCym
F4roXWH84Tz3dmRhysUJnrXgiiGC+lKx9AFDiOmyFfBMMS/Wx5JpfCp7FCPOxutIos/45cRolcZ7
T2r2A+MVW7Rie6TdQZ6/Nwpb1Jq1mdPklLvQ2VPPgdVczNItZcJiNVMudSAdacqZVa6yPzjWHpTp
EE8aA3cPirbcNULGTpxJitM5oFwgl5W3K8lsPFgxVZPH5hOS2jZALLb700LCgxcRcpasxvOBamR2
AX/T+y5Al/wUwyVgu4Sw4WqWeDPAPHNskMQUimJPj2SL6oOPRZUV8gIovEmjuET4OQbrOMwXN5CF
VopGyKqCtSXgy9tJRbLkedYeN7Th1+Rl51UPHtGDEnAfa6uVlnKCyx+6XJJ0qbGRb8uav+fvZ41p
xTZ6+fTg/foZbethPF6HFNxJRMxB8L09nDTnF6NQZzjMqGhIG3gA+5tl8pqv64RuX+LWXeNhhuce
tBQGJUhYHrokFEg7zQc53AKQKEHhKOrRbiIMI/AL+hP7V5hNN+0M09qJyS7oPPXGyLCrrEc6uk4m
ENUapn3Q6cctmh2QCTYJUgkQmkBoqXQGBLlIzhQMj9cx62QExfHE1emIHKzGoIqQmdpGXygUqJyX
4gZ224StVTwZ1QB4tDY/yvdWKFr0cLEcx4m5XgZguAraGUinpcR7M/NG7NRDpp+hkFB7lYAbyKN6
xDCzGn9CnkvPjDHU4ytcLxJR1eWZdNrT17Mg8THZyW2zVJESXkt5IXQekYH2YgabcoBrSERQni3e
fkezkLjBqu4qlgCNCCEFgQfcfsUNQwt2bsNinS+sVoRdiM7RRAFl4h5iwL/LVKWDTur5pPn8YU+w
qizqFHz1RKhCRZqC2sDy1gjyqSSgQ31pWKBCkOz1lMpEX0GlnoWFnDwdo6O9H7uOvX8cX/akGbxs
eNnafmd/iQZ16ueZ3apXd9poACbVfsKoe/KxRxIq2jbaKs97n1NA7hnG+QzVGRnPrK6iDVq/9tlh
pdsiKuIy5KB5+cX8bGbIYT+uR2DVvNR2H8PFysjzxK3vjomj1ZZURUSE59vB6Cy0Sk38KAK4646t
TwP0Lg2zhc78MTQxSSrtxbLvmJQX7/92Fll5Hw77rLiFA24KThCJmKIgctBbYwQu70cOv920JuDR
omxfcOuYjZoreG1mY6gTH8FnJXzlnthnbrlTfo3y7qJGD+rM+t7/hDrbDpyZzSrIK+03gDxp72fo
OwZcVzHr8HFVauJlRtkOMgx0yLzqG31R6nuDODxOjrvv/VhjCaj3bPiGBEksJSB4NYZDWf5kZeeQ
Wd2snWe52lzjIMlHYcJZKObMXY5G5di7x3Ih63EG69SdoDMRVyZHaTP+/jX02f6RXvAxXi/DyKXi
v2I+OH+M82kgyP7uooh13gmS3N9mco/jD8lkUxLAqYtCXWncp5biVqyDerha56jqvAVqfxlVFsVa
t4EvWS/wh4xhLIME/dS+UgG0btbJWNvo6S+4Kj1beGnGIayyNwz5P9xsuZI91LKOLk9+YCm8qAl4
MMqH/zCWnWHWnM+pWV6x0nkrL5POeoPIqLrFCnsYxXXkuhTSZDPOv/nbvDx6Np1rpk9WBT0aMDdR
IX2UvMuTK0vWPDAh6JvEJddMNMF/cqK9ebPKbuoxcJBbp2nHSmviGG9Uz2y692zWuzFnZY4yUYbM
75+kNClVkVgm3cdGtaB3YXXdRgMC+DLUuSPtPh5E+PQImWM+9poLoqpThxmvYJr16p53KVH5tr+Q
TVP/4oZ/TPtMUpFRUFrDfBdN3V/ZmlTw4W/t9zGq/i8MdlUT4c5vSIyq7A2NA08+7WLnR2KJqNKH
Y/w/+5sLy9vaczzn+t6QhLE7sgDfrdUroAGB7L87le0/3GoSsA4adgwfUQnwUfuIlsBBydM7HnZz
EG9OQNFsVsm29VwTrPDE9yZiKb7UFzm02kzQxjPhmZLb2J0OMHilEnADL63B2Z6pcNtodpNByD2Z
EZdsVwVSlaWA98CdNKdC7YuuC8MVxFUJCw6U3KBZtMPyLTbOADS2kD7vXUc9ngP2j3AsSW0rcd6u
W7Sr0pQnGnwt4fUmPFJMPLZX7kWikWME0a/GZUVKiVPndoRysiVGu+n3KL61UjLAgIY50+pkFPwu
Llz+qcpNoDk8ZIqrXu9n9HJ5IrwGC2CFb3J9re18x2etMdkBlaND6/Qd2fZu3wmzUc0x2ZFeuLgq
fsd0aNCYAIdvAWwYLoizCtX9U1/rbz112UU/uG2O1wLhoH2d6LdiHZrC+r0w9vvUW7D3BQFjOoGX
I6TmaVeD+DwlhGL14bsD+xneJKrEhGUsMxHz0oFpT24mJnNHLMbh9fDyfoNQRsnRMVEpGKd6WMUN
wD+PdIgEgDoPZ62m3NsGvHdhXv+1GRkBOXi2a8Hs+IYpSMZXZQHY0WrqIyQdCJEmuJ3DiXKcf4ub
33vTEV8ffQiofYoSfsJppg3ZJYzn07WJGIo81jLmPdJxP4XJuXQTFKC+alSuNch45YuU2f6JoSvV
zd3BJH22QjDYoD3L5Mmgku6vT00bRGJUXet3sNbbzeUnm1lGvMKxr8uJsrtrq8s9yAVkS4zpO9DF
2tXPBlvEcP1rZCy/GxnHHlaFNRLYEBmFyG07c4n0oQ+o19eXUkzeEgDdHfhnWvRUBHbdUfXnaxGF
8H0WrrI9v+fBqvIZU2LJCFNW4OkiV1ISAU4Q/fj+4YjpUKoYbiLFT3XZqRKs4RQpW5Hi7acjD7+4
O64X02kdnOqiSBIATTRcWElbmd14ju66r7gegWAzGukLjZv6DI8cMEjGDhpOby/NfW/YxXZNOfOp
22fpD7QCLDu3KV/Su7Z87WIe9TK2MuwAR9gcqzF6uAH7q4/xdy/F/EJgNB+pnKXBY+R2caKXLD/+
jcLqwxPhugq/eb21izsGHX7+eEO0RUndnm6yFYi0ls4cxX7oKkAaXiqPAiW5kI74wRn5eLsshLBx
1qf9/WAgP3/z+fBTDuEooCcet1MLWEwzYMQYPC/Pyx49TqbjF/ocy2zXyUCER1G14yWq/7t7CWn6
iJ7ebjKG+NUKOI0BURDvK55n8beU2pWQslN/KYgH0lKM//4cRvUwzzIfQeOIWnpOarPYaX4iDyGv
a12u8VyD6vbvW9sjH8Nt9CDKEW+zDu4iGcVHQQir1qdmG9aBu5gPnQXvJED1V/Ft+tj5ESCtUcJN
7d0LzjekSx6vkDMVm+HrGDMjtN/02uEe3iWBuogSAP+lMpn4aK7obEw1yWfulz1l5/JNlMKbFyYl
x4scoMDGLmB86CJHn2pTrNCs20zL2hpRKBIAHMLe07zI0DfE4gHr+FS4xj8bGozSluzLvE1RjNr9
69nUBEwVQhavw6n4J3CGAAh2De2g5hBWFJ4atTIsD3A5shXreOmv1Vc8y5kV19/GUnqePqZZmAJ4
PrATDPEQdJAZxZ1SIud/YgRkLAVdBTk8pm3EuE14ifs9dGYnPmBvllhUkaCFVLIzALZDbV4/sib3
pi0I1BJ/eQ54+SHLkYIcJHaUoBYX8mW8cULvb7mESoiciMLffOrYyngWg2stbie2ooE4yJOtxQgo
q0xH4jXVYyAbzH5FaKn9sSiJ1+yiHeRt2E86FeuC1PMKS4zDIKexvicvOVvL5FEPtrToVvYSvnvF
FS8ivUxXUL/r9AWGiAedOx1U0nA6lU6cTc7spOvYFWXR5H+hysD4GwYq2TszZpt9tVBrdog6PH46
qvVzLGB8i5DGgKRew0cNsJ+/c7U6E73GmDKXtTQFfBEbopV+wgGpt6eQLYnOjglsZ9qIJiVW7osb
8gvfiP7Iiihx7UU6DQCzqKajn9eXJHgSS2/sYWkHmE1QuS5Z4jQvPLDYvzN67vnNeXDbtHlHL9KK
qEpHh3qn7+aKytnt8zhbdwU2y+UpK/keQ2EhI7rtlGvh4Y4dqvEg4FBlppMT5kMgsP97DuJCGw4O
6WMY0sXwRWseLsLYhwNYG1GNb70AMOOeJ7lwV0TPHF3rITH0y4ukEtLVD/78yzvedWjtwPTmRQ9M
YNv9rnng58WFpVODx+WkdcIe0zjwfXz5EuVDZlE3Upncwpk/a8XkOP+3tFlkQbJ99AsLL19rAhOu
2TSqgXbdPmHFxgmLoWs0PNG+O8KPKJvET6A7aloI487thN/vjUgn8wk+XDUrh401FAVPDtqut09a
pGxzyjanl+RJV5BFjRbPVBB8I5lrWZHkBuI6dLQzwTO6l6LVNDZILtUYDbN9YoGQ3+I0Le+TWrm9
2lnuCWQOMD0ZNHBBezju7Xhtas7DgaWGNigC3CogENANvzklxnVSK0WDfm6Mw1QLlDSwcsxHY+5G
zH8dd1P9uEoQi9USUQ0eYqgSvlON/j57KipBJ2cVIbVo7dx2tlHexFEHM4KpLmA+4dPoXBneo4hZ
QGeTym0bwgPgjRAKwmF7HQCq0NXyfRTwU3GJfN+y0utc4Mh4Pcvz/cTFZEDfTKHLt7f5YW/IqqRH
SaPIO9nrHEUbT/keNJGI1VEbMjsJUlu1NZ+0KlMVdxCX0rLBXrnFH79wI/7PcOYVREEEgRdSXTTg
BdzI3yZ2JgK4oVUOprYHWW5b+7IgkR8kecbi5uq98tEP73QyySJ6n1fO6hOWnpm74mviqI6SlNnC
6APVp9YqXZM34pmdKQbqcEF92LKffcMbLDuFMSyWy7fk8ZZv71CJSUweuVbp0tWc5Kc+75F7IZMg
n2c8TavhqZH+7bZ2CRzP12yiLwzBFOqH6ccVukrchacIwURxlxPF+qFYXYSp6UMHjUwCKXr462Xj
RzCm6yFPKUBtxAcjyWwlD/TxUZR4zSvbPNCSKoyC7KSXL3YJk9saOwIqSxFxva+uUtdHw7ikWnp/
LHMPRKV4RHJ27oAHyJl6bZDX95FGgJMwDQHVpZG2U9JVkRbdkOxpOI1g05hfVdb5l7FfCWc++auf
VeORuVD/yTDvm6equjH5/QBBIN4M8ZbBLLxQQbCITEQxRogs5i/MPR/lD/tsWnZDpdj6hdeqOaLx
GiXlpsFol+Efc8pRzPm8nDFTPP7wMvfScdPJ3m0t5GGe4kfdRY5Knxxbn6S7FFwtRGgd5o+s6B53
iwTdmjRJwe9JfQ6fciMQ2PmSExj5t0krOoAjd5wtXNH6KKBKIN5nHsEGeFSwcN2vqtDHaCXsnN+V
faQTk+K+mhGhpOI2x/KERfB/nO5AWIbcAwUGGfGlTkpcudkyJPkFv0coMIkU6RjwCjoL31d0e66s
cNcgUJnWVM+SXbLXYLOOzh2KNPZdwGzodjlZf0/pmj59b5oHqpH4VzwGMDBOFwnp8skBHSLyg3xl
nex0zGYWBEFYqC6476bS1T5MnHwd6fxjS/LH7X1H+ejFKo0dyMi7eWP+nsAIQu0HGxo6TrcfwssQ
bLvnMxhBVGVIPAn6tlG8r23sw87uMwyU4Ed+oidPRCZAqM3IwkmoVn0zwKaT+p/V9m6BjtUzzVdw
UEd4Irx/qobQZtUF0SKdQti1zTNyk58HA6G3jMZUNiKHK8KGI0pHabbSdfrzGbz2igYY7L2NuG1/
orpumFYBJfMwm/Jy892mpQmdFwPEywi36c9o6bvR/98xxyDSLoCNMigq+F1jsg9yZbXUoyaLSO2N
Jti+aX2GBLjpTulhEgE4twJFca0DOmjF5q7nT2Xt41TGIC3mncoKoDEC+K6JKWTdFEwm9paCOTj6
0N/xRvOsH6ttfXrZxJGrLF6+Jl13l9yAY12bxchKKcXscYVEeyv+h3v3NRe/0RbhvqWn/b/hLT/G
uwdy1AWyjjvC0hinGY6REBqZvvDEFMA8DhpizeHxtaXRbUOJCkKQLO1o8QJvpC0EgpuckiXh1Lmd
UlL5Nb7mNLFj6B+4hkzqYWKorq8f7Jp2YLbpN67UElygq+F5LgAfLmw4z44DUwzwdSKTxA+dpTJj
haawEwxgkpdS33oGEnhs7e0WrPXLyXrMZ90A/Y1bJOs+3Ux1NaSCbtlxDFMUKtB/bJmfMR4UsLcF
0Ja5E24gdQp2uZgyTt/zElph9rKMKQDI6OQifpj19bnkZ/3TmCBuqjTpVX4xRxjAUWYpnyOWq/YV
sj71Xc2vZde1+YdrTQ8OiwB7041Eyet5Q1qBYdfWlViEMEbU51HCSkBfUmxa9k1nV4WxaIexqX4W
ok0hYK1ppta9T2bpOhmEhg/7i6nhTUpzEML7MidmW0vlMEp56wcdLicOtX6b3kb/niaX4i/q6knI
96IxB98QrNtpqKLz9W80Lx3xG/GvvzJEeT8FUBO7Gxy6yc+GjvPJQRNur8ldmoOE47x6ypTxpcX8
r7gLs30LBVhYMkfo2biVvPC0KKt6sGKyQbuyV08Eh+RMhqs2yWO+sQNWfmK1Rxk9MHs4jj4Mwa6x
7wvbaLZsCiaQ3rXY4VJkybk7Y7rWO0iSATfAyYQReYqbGxQqsDlIswmB9SHTn7tNzFrVRLQ4ksV4
yo+w7CR41ETnuk4EEkEU0945k78nx2x3CBLuLMig/JOYEh6IfIqe1CFwsFPY62Y+o3rpYsc8/o6I
7AvA3pn/IdMlqrFPlm8Jjii4W7vwPIuBjabgAvS4uZ3eTxBd50Orr47jju3WjiXId73K0vtjCqQn
gqSOiT6QwxQopGi2o1UO1/i36CWIAExhhv86CTtZAFs6MLJ+jbfjGBfSxfzQXAn1kGc/U4I/GvRe
mbZkCjytdIzpxWnBuzmC9j2OX3YAQY2ob+iUxQeLMv9w0BbR/puIImO4p2sDFp8nKc+7Y39apFTc
MBKP4iUO0ssR0kNKrHaDrEKhZy+tmKR/eOE+fX47SOz3xPvUTqb5b35Y5UiOX6SjkHFpCvIrqhOA
D93lNlDKHqNviBTvjSP7ynUJc8Ks+uSZLag97whwk0AQB0TsYY8U+qVU7y/T4Iq9JintxQLsXBVQ
O5LnYJXtAV0cOfRMGTZ9CXNkz1VP3yYTY82qztZLkw2dAg5W/lV5tRNEcS8wa4K0LuJgimqzqiVv
sSfxT6laBBQuz6/7Ebh9Ck0q2+KxNKaa9CLtj+DSCitqDqeMe6/UpvvKcjihSbnp0nKBYQ3D/5yD
zXbdFr8rEqV5/k2TYZ/WJ70kW9HwqohSfrLVcPcboWmhjzm7XV0+7LIgTLAt58vijabGgO41YeNF
9whmCnKyHOP3g7cIKyoa3AnjZDIzoWG6jvoZTdIPvDUeaiKv638MkQ5qaJDTb6HA7l6q4y2co5zt
u25iNtVv451AK6oQmQucX+wAMf+NPdSW6kzHLkzlKWyUetfBNwhaZwBoSRKzWh+38MJUo7juLCRB
Exh9OUrHL1HaK76w9AlHpLSHvGpJkl4r9eCtKDwz/oVQ+ezAkMLvsbhIu4aC4HDn/XtN3uQEi0aF
gDUcN1GfQDsSmy+r9viqQnvSWYX2dKHBRV9Lw0ErIvEbaS1IsvFhui6kQv1WVOPil5qMya09UWDo
C7MamZqaEWhGzrC4b24sxxvX8OhH+nLO2a7SGu3a0c1G1unzNp7WdSCqROVX0KudVMemBJwX/sEy
X8b/VIlo8jNH0fj+QM61VFrglS2IJYLp3vzxtgCThXVGIZtbnTR+33ffOE0abyBlVhoh1ab1XXLT
CMbLxcwaKIlYrVSfeCZ4dm/wr3AvvX185eEOPPB1nnlqHDdsf1JM6sMJEaPdX1QtU1viZpdtiPmC
KUmGVmxmOTy/AG7kPANgv2laYQwfry38fkWaD9OaQJvz5qEs6+EvU4v4om057nX5yN5rsmWtRtPT
bGt3eD1MWXsNXyEqI1V+YywXD1Q8rv3lvZy1JSK5u6nAZ11AYZgNrO01WsBdYtQOwCHmlhD0s2b5
1edr+j6rmMx87HjkBfUr9shF0fgeWmhSq7xGhCKtgkpcYUxV9olQu8lt525PFpbWmH5yfOAs/Czi
CJJe8V7hHc5mz47maSUdY1AjO90urcS6s8X4iUf5EzDLEh4mBZYZkM0sM8Y0ZycwtqBevP6xKJ+l
gbl8cx2FMNnNlbqhenBEL7fqiX10YTm0e4NWl2ulBKin5SAzsleiOifQ82PEGonSAsdiNaRc/IMK
+80mUAIZSNY2hFWEFfjLEwEvXGGKGZbYJ6k8qHyyaU70mw64FUXc+vcNttF/MCJrZmJSXtRKDvjW
9nJq43NS568+ADznoQkXELuutIfs+naUFfaZ2MA7YIak/tYmHJoI75mnOTokkL3Ntzo9oO8xunSA
iUdQlvKENKnPjyx6Y1WBg3Hra50ak6Vj7YfqESTe2Un2iPIq3S7/SFWXVnsC0ygaqmB29gA7BmJr
PSV8C7IX3Feym5dt6Oo04w/sG6SVGzelgBCcqHVcpkjTs5LTxcyevIYXv78PfUhEUySTo0mU/zqD
7R4iffN0SPXlX8VVjs3mFLEGbsc4FPcQXq2NM6zL7q0RGnfETX1FwDTQ1nrbX/8FC1HJrWDQnxn0
aKFLxFzDBnC2Go7Zs+91S2eI5xAbmtGHLAOej+CAKm+Kd7gfLTdywsAN0L8svqUCjbyWIwLJZK1a
qUjpqYixlsXJ2ZLkZV5a9mIAFfI+DPm8puFKaRJnALpVcIm8LxnMFTf7RKA9yxEmqIVi6Nxxf9ZZ
4CZyTjTk23Dcwvb91jNerzpQHLxhMFY+UQ4CFlPeeE8O2f2SvRBrfagJ6BcpDGAblP4QAneKftTC
ox2+Tlk73ZT2bZ9ulPajAqgTv9UB5l8I7xnRzHJh0KWcqriNVZhKAGh536eCuKn9hJJDBzXVx5f4
aabG0/YTC6ylXQfD1w6rQ2QL0ikN5Up6QOVZP0F6+vv36wuc+Y3CkdPDdloEYoNc7jq529Bm+BA6
m8HyKL+H26izrwRfoeKP5QVlz7JR+dGFdoM8JOoBB0x8WDrjAjmUItmnmMlVaR+Ls0OWtRCJEGCa
JIe7ZaFSnuBH9cVsC5E3Js81J00FTjc84pGCwLidZ7MbxJjP1cPh81zcVndkRAoFWYgGRdgrBRXq
Eji43/oKHp5hin0PEsDgVxe4aec/3BPH954ceFiNrrSL9ABN5uKkyQrgBu47v5Kl4FG86AfHDeM2
06FH83zapipxSqGxr2rHiIY8JNTPfiW3WVlWKjW3Wh3+gLY3JJUsY8NXBjUZNdNAotbetWZEtyVF
OWjIfHFSMpoJCH4zAU37bzvglznPqz73tKLiahCCRrgIlUAo7Z4Vst2pFYfxyHQR3NgYbTN58qOd
5SEtVTKrcDqI7ppQP0eUxd91xJouNW8Fr87Ng5bSzDTN7Z+PScv1Vy6HZPRkffjBiuYs0C3vWfWB
K8IvZlXBghItz/0j1RsS6mkIIFVoNFE5mGrIBwK9EeLCAGGT8hKSfP7aXa5LYP6HcmMmacTJSWsp
3yCezihRWdwb7Apbx+S/jBrtKsLnky0oVJ//csS1OTeCLhiCvFYBoyy1Q+AO+eAA1DrIlfEzZAyG
hQMr8FqWzsNDCmoMRD8vy1UwvsIc7BVl07wehG9SrCnhzdDVmRr2uKZ7+F9g6+ibsKcG5lebL7YN
kunYUb4+dBizgbHK4CD0SiT6KX5vHr1VKoHj8C2vUXYxnK4NR32DMFwXDpCWmcx5LCLIT7xQWh/B
ipio3nbnh1Kp0qYql4mSN9/zsE1YgjyanKmt3ff57mMRmm+mOiNoDOBxBWRcjA3iKHYDV/rDH/NR
GpVjzsdYUbmCd9/fluAF2vmA5lGbSb0qxhK/uMFC2MNSDZp1QVjp/HiDoTkF135g4gLIpLavV4Sj
AZ/bONldmTyXwXSRPtNKqKUd3mYNY5bpyxyADm3DddG4rXAQWaaQiBlZJUP7Q2LsciVtiI1AX4AR
N0JD796Gox6ECRFqlFSCOJw6qfr/1BC/udOz1hiTmOYXH60LdD9p+6XGw00ANWbtOfEoVUd7CYl3
kwoX8x8LQ3DeWw5bSlKPEGhX7RyEtZY0+HWyxsBeRAv0DE0D5Fzjq2a1+Q/DlL4MbfQfuHDOXfLq
2zyp1KpEqMDk7tE7o0W8Pohi+ZoPf4218daJZ3/yDGa741r/CDxUCZPVBqlQsjZkBCWm/T7IHPOp
aOfCXrxubnWXzm4PQMnYFbeDkYiooXwLx7M3+Zqy3N4I0ZiqfumFj5m03pkn4JsXPvF/5UtdoPsT
qOihyFYfGJSvGrtsIHiFtXxoHrenfqD81o+K5WWU3wzHgeHt5iFsM4FyXnkeoh49Zn3Nk4GDZ6P7
U6Qa7hObPdAsKu8DyBS6J5cCxyZZ4KYM2ogZfgVJ9JcA/7dLfGUMmphYBreGJt2k/vIYgwW2idiA
TE5DO+WRCQRBqusnN80cIqfcBNv+g+ytAs9CiIGltBgYV4pwu/EVh+NRpTBOH+tk2/nLSdc/t5wA
s1M1V5a3d9wdvhjNyJ8neVa9fdM0AS2HMyuqULbGs1s3iDnPDIgtbLh7Yg8iur8iyx7WdWcnyev4
XLD4qBhmjpoCo6QdIKk8g5wM0SLkX3gsU/tL+ht+R+iM1tOtMtJH5HkstEKqCof6e0/PVmKzW9Ly
MxfACoIj0Fwr8jIgzkTdrLYM8BQ4sFn4uiBEUtQg/YPOS87k1y8+Q7lSGDuA3TtYZS+GI617f/Nw
V9tPqSyUc5Pz5jetv2OCnMH9UI6f8ZHR6rjYUq1Mkp6QhjMzSVBUiqnQ7wvnzaPRCieWRSzkKl35
UwhaCwufkISKfHweY3dAcfK3RKUg5vgNe7SktSdIflKh0YYKkJcdTApkHkcbce09UiCL3s6QKJlp
580BWUfELpGoG2XHH1Xfkx5xN+74NtOkbowXHJ9TB7p0xVCqdsYXNgKRiswZIWPpwYH8LzUj478T
x1TfsY7HfIu/lwQOxaUtwbg7KimM8LTECNTHmr4oF0H5K5J0VEg/+d1ydJa3BtF8oBHv3PiGfm/9
HawEa53WQ7w3JHfY6TY9WyOAgJnlaak73zOG+GXolsJ6YA/ypJzlv3M/LMzi5ACdXZSsRP81Q9Dm
esMNHYoo03q6etEJUt0+RvPVpyyfh8D9c9dAG8TdQU6jbUIb+4XzhPDNN5XwQe/1VVhqZcNOIBQe
wZw7Cxi4FiBcYJ8DpAR37zVEYQ7xKJDWuI+/B3re59hJKtDvL6JTICWVGdgCTec2x1ZD1SQhQvNM
xwsQMeGPEdhgLpKt2UCD/Gcu1AzR3yaZLGAnuE7WuBL/M6r54OYNYZmXG9NVX0COp7JDXRplNYW2
yYOsZ+UP7+0S7uTNF3iRShvgM7rJ09V6RKItKT3tYXwfqcnpJsW9332hbIOnGFUhMVSBSJSxqKP5
+hRcH3R+XHmBvZnr8y9gj1CBd8Y6XCw7dOEJvrYIVQoqiS9TbqdelH/U4q2Z6Af2xO0fqcUY17UL
b5ZAU1qmxxUlP5kWn7OJDonuofamU/24cPEOMNO41EVB+j13j4t7BYo/WPMdOkiQIuro8j53Q9Ua
phFoOCDLgV5Yw3fWFhsFMyFOeW9MZ2FXgTUZwIJy6tDsFB+oWuzKzDX75IudYf3F35KLEDkvYeHx
Hp5MA2rS97QPlcTz9MqQQ8pmoQ4VfoWnvwiLKO9NaGLTihZJ9ad95rofJXPdcfVFmfVHryM1lOL+
Uti3EBcpzUJwLcco8IV/z5L7j1yNfR2x/r4Ep06rZKqAI9QyRAjl8PliOSspp4470hAZxewZ4FGX
iE+PAPQzxly5gddgbqPMLr+X50JJ8GIC9ildKAOcdXN3TmDZZWyhZ9UWVGGOmcTD1IlpjpZNKXXc
4K77aqkK4iSBzhK/MC6rDmzrsk1PUWZvICSFBoe0A2TNvbUG0ITSLkcIJUQNNeyRoNjf/EiK1J/n
+zhfqDko0S/GAB3dZgglD2bwvHDkz4sr1++CIv5dib/PsW5MgfiYzCWSdHmHSzntVhsRO3hH6Rd/
ZlXGAUge14nhKvKMUPjiRBq3NpPa+nU54rSJM5C0GNHIqELolaVtThYeVRL6LaQzTMc0n1ByUAUK
qdZIHACHB96kTq+dkcei25KcQS9tRqjlU9dvVFNnOPj0OQRPZwC5iyb1avO0IUZJdZ2fRCez1pVY
r9oSaI/0fwpGJL0mPEl+KVxg5qw9KyMH9GdgPwRAfY5YE/A5HkhNT7mZj/oYS6fUTYMadZXRJsJa
/k+5nOyixbZOb3MVaaz9zFoqoDpzYuT+lUoqN1G0X9SYuyU+LK0L9L6yvnAcXdoDQMn4Mv9+8RtZ
jnxUdaaXQrRhEP6Tmos6yxcKV7Ez6X50pfLKGCAeGk47/yu0q2/LtXRm6RTMlQfwTWJTENLl5KRu
ihdjqfd+FiwSaihR7WzVke5sk57thhNfakwi62ZdB+ycRue7XI6maqy1V660MP6iCRcrQyCmUeyd
S4uw90WlXf5z+Yv+TmJ4eH79k1gbNlLfn95gMq9Rl2HVMUA5jBq57PNANpoB9rj7700m3sz42Y9s
ZO/pQTRE/s6oNkOW4Kn9+IHmIvlQOvCfHXGhRVIHisjibDcOgeIheKa9rfOS/eaCbKSIwOsNrxnw
DZOHyCZscim37eo+m7CSbg75ggUHkkWBEGzqx6eMa6JpI8ploiEKKgovoqF56/qzCT1HS10hWqg8
P0b6ydKNeViW1MdrrVaoAyEdz+K4D4tKk0B8lFHpJZZVyu7s+/9ad//U4lqTBelRAz/ZEwb96NGr
g8WyrcnPPfNZipxVrLAEC2PzyekuCsXZahaWVQumtmgTtC7j2Ol+JwcQqrV9QbPiRKyvZpr/bBJu
BCnCaVBZFlIITxUO45zIaLkeiOFEc9v4vt6OSOHrxc5poO7f0uyMPeHU14B4S6jH6P+xMLGoI1jk
r8LYT/EljecB4Mz00xRR5Gxwv//rOf7popYxDmauJHJgj8APdTlxBVAzx3Z5xIFMhl5HgmwpMQRe
2LbsR/0AgfWINoN8pKuFHItLykbJPdWtzOM7crf7qIIp2RhGFhJUXU2JL1qHyrJdJCSXB2FmCru0
RqspidGYq/o8MS8X7+L91gFSPCzEol7uA8B265sjaZM8+xJ+pwtRaK1JmWeTjPZi6qsbOtBhgiIz
QhIsanqtChGLewQyTSz1ILy2D/6dDflLU3glTKyDxdx0WpWD/sh9Pw8aVlZjMqLWwQuq1yREigQK
2yzT8NZ/FhfVpU+9IDW4ZreeKWJfRgNTYJygy3tAWJclcEvhb76wDzZPjYAPg0xYDRewP+Jn57Pw
OxgTSJZRnomyWjDsLoWr5ZM6/a0sDcoqLmwnFArUq8eSCsmQybq+M5mKW2hlWp1S+6vRsp9NroPO
pYX7NY93GhUWmB1E2TuPASFQFmSqiJ8xgy8HRB5K6rhB1pb/jHe+V1hqevx1IfuslT7Tn6f/sHCZ
pyYhAMQ/ODgoyDfGP/Ab5GsTzRAaQJD4m9VvuZ95YQuZT7pplKqde8grrMmvNkVcrBGEhhBnC5GF
i2Ebkt6X7jhweseTR1ur4DfSAdMfTzVSJ5rEEMFwlkLGfq5Zl7/SLM7/fgDH3NnRI+82yMJTO8iF
a4Q7RpLEeBAc5Mw0exyaLSr2kJFXf+/llOH3iNPe20XgUm42i0zNjFirZCHq6IzDuahJoj4wZ33D
ccAz7hXGXQ6h3zvP5zV3ydX81rW3wlXgx9PlOmmOYb+UdfRFgcPUm0ZP8dWO/zRk2wyQq9eIGUcE
2/ccdHBkOg5NR3mxWNjB6+lnQUdD5eQh7nVEklJ1UvD72JmOcEvtAE4avKwRpBVOratkRWmWaOIU
tHIDOS1Wpx2y/dmp+ERLk2UK77n1tbg7K7stQJha/cDSy33cm4VED+SlZBkTxPmWF0FtXFezVIVk
Iap+hN8imUsGWhEDROMSyKOVnVVedhXv5AW66y4coZjDPfKbbWgA7Sz+FHX99Z0qn68Tz3M/3nF4
8fU0b1ZZ2fH/2ZR89l2kfbM20Me+4AFC8kZabBnvpsACumFdPNjOADB3ZNTyMNcSnxSDw7UhpAkV
f6bruOqOJgRymaAYAir5VYrJkHSprUCkIIyzL2anL37ZuTSmFOJZ01CNJH3ZQ1lXIvEikdFp5RVt
7+ofWhyYx/4ivt89wOO41Gtpicxm9Sjqla+aP8fqU2QuOml89xi1zJQcF6OoshtR+BVPJvlqarq7
doe/wJEdbQMjghCyArxXogeAfodpvbUzsvVvdIPU9+erdC5/s6h5xrAnYkE2Hoycu2aog67ZSAe/
9Sn+FE1ZTH6eAGkp+RJfKUijr/PHH27Xo7+BPWxM/89eE+n3vNqGkwbOb86E4UUY2jsl5N69Bdqh
iltrPJHl7p4oYax2Nso1Hss9VZmJSXZ1ExgSruI5Bv027xrhTK+POzvvugKeELqz6a8WyJS39m6T
nYYxP8cSNHfay3EJs7Jx2TD0/RhFc1E+nVa9CONQzuMGQAXEa7WP5Vaj3ZI2ic4nOLweoHPgZbCb
UHUppO/NcmflkMmET6sb6LBwz7hi2DalV+sYGEGHBc/lVvejiv2903kvYaPLs9zol2IuyuG7cTZ6
UsmjCIksyMH7hPtsQ3urUxmP+/g80xn5ENhk0AisEj3m9EBSrc67or6Bv3z0QN5CkyGg5S8x77Hs
ktbpGY+EpOyA64xH/bWbesC/eJuN4k3Ijh7tt0/2e+hKtfadIbK7pyn0sJgDYTgOxGAlizXO24ue
G9zqicu10wtoELgM8P0uc9f4iPjd0wPbllfSBG7o+7Z/ttVzuWwM7h0XBbYENss+QCp49x7ISohl
dXgJeK582PskTrbRGa73pkG0N81o09RkN+8t0tK4qlitF58rvbd9eqcdq06FushCQsLRlFVWzOWv
lZqA43QxjXOyXoj+DF33JKjnWqQ5VC5kDiPN1p/MvZ6oFK64ToQ7EeuGqAgKAhqkuRwwbx9tM0gs
vTr4AJdV124elmVqsFF7qWYNu2Q4VaMWxmFNFmgLwr6C/8TPckvbs6qEz7ChLYjyyTj2jUEXQsZ7
afMJrk6mjuOKYQ2NvRb0NPb3FZKHAk2N6oqVvMH6JqjIFuEuLitxvmaCWx3mcP2oWqrExqF9MP3P
kZNIeitVv4X5VO0dW+tMAtMM41v6djYT/7cJo+L3gcnt9cRIUuv1SXE4Yh/2FhBV5Eqo+/CHmh1o
cROJC8PM0p38daSeZEXgqz3mWzyQ8IiUkGSXRwMEBz5CgUagzEdKxSwZeP6P4YWvI/kcib9uzLVs
11+IGw1THSjzvXkzyd1aXSOIvdoNH9pzt3yzbE6wrvLnjFtQzrXZizIeBbyeo29Mht0gjgeyACuh
XsQuWsxQ4KQInzvNZ23aZmY1SAr3P1OzlnckM1P3VViO/UNEIYztCzMX9zExd+1/wT/cs9SQd0mR
ErkEO9ZI7nuHERT7vGCyAzWQSXW6Dkmxz9SPi45Y9sW5J1toBy8+O65iqIGGK9Ebzp5m394QGhSC
7AxDVRcPIkTCr+BJr4p56PISAcjkFM9LH4/aZ5vy4rDcP8lCuwcTfCrYUrnIuH4mooAF7pVlsoLF
Sasd0q/CCRSYLAlrW9yOgUqrlg+rLJkXdK09OGETBXduCfFi3dkI8hs/WlNUfzYcHeeXeZwQ8YAy
PAwnFiLBqzkWlGp6vsVn+6wo71fq+4g+21rKZagpLD9WsZzWwwMAjwNHiDf4Cimfqsnva7xFsuku
1yDkmpOiLfXhAmtJMlUtaeCOnSZSzuLv5cS87peGSx5AWhh6d8LizU9rDdKbFX1dHWPFJ7qFq69R
yUTCXZA4VRlgxopsQfjPB4XjTncG6TGgzChIFUaKpz7ZftKdsWp888iqxEQ6lsfpVeHmDwQ4XOJQ
DNwLoDGf20jMgGCXIrv+newpMaUTNJ2DyEAgOtWI9Ye4ltUH/tq0BJegARmjCoYrvUhnzmYhwFXe
+rw5+cRqkVDCBZeq59SY3aTxxJ+j7PIIFt+w/ynyrbiQNUqc13FcaiKhgx1Od6OKrpmMhXw4UuMY
qMFlKR1ifJwsnIyMbBn5uQob2EsTyqBPORCAssflkQRZYgkFb57ANv34DM5QY35u+JMHCUw7nicd
Lx3IXTNewIMjLarMqG+F00EGgUbQ+ya2zvU3qKSUsucyFYJF4a7OXEH0fJR/dBeyL8ETTdmk+kWK
ZQjzXHk150QEonez+pSNa5ajDcC/fahJxWrEjm9sMGLAeYlHGca/IhZwZD+E0twSMtyggnGaPr7+
vBNoz8U19UeafD8hK6X4meS7CNP2M/l/29Goa/z4nRQ6zsZrxCodaU3km6LwanO0iDRiwL0jzZBC
TFaa+S5/ap0bsjKCjKMqLYenZcleV8uEZzDSekDjWPPyWs56rRFSpxZkW7a0cCCdLkkUaxN1QUr7
z9JC7YNlAbqVbKTmYFdJVSS4ziCG26cuiacDjTezCuEHU+2xilsIkl8hd2q1xJfNdQlf3TgpLceo
AllhCBRJGX1Fuu9x8luchewlYsqFLDBB9wleTiBvfQxLmDrROmShS04bWM0gu3sfbNcrbuw8aDc2
g5hGumvF4zIkIM3xc/a3HYy/smT3/kF3VoUQV5aa/r9x+32E7/YqdCd4qJH4xTFathsH/N4ZB0Cu
muRbKMV5fgl4zoq0XR2OsHnGscUA+zbwIHsIkdQVvA6QYE+jrFtYVRTkSxeiYogjfW/PZg5sgG2m
eaNRWxEsd7v+iXF20b4IVyFy8T8e0a6YXTtI19kpCv3JIkF73MuBmKZY3TwIFOJ63cOndmfFjx6/
ywKLdjjekoCEWEf8GLDaMWv4lmDXgvaHy21YsqGD99YL1CwIJZsacFh3xLwW/Cwvu5pB/cdFg8dP
bh4TI0hRBYjNVipPXm887Ck4eo9qPOVHCUHLNMRavts6dCDtLVqfrG9bkfrxfOiF0tHhlHMkau+n
aEIeCc7gNpawsT1S8ib/KhdeJ96YgIkTgCV0W9arADBpK56uRo8ktKkYD/6DPcLrdhBDyvtIFzh2
tkPkKNBt/b8OrpZD3Mt8waZonSk1KFbDCSPA9Xqn1Dl8DNxhYuFhqbW/GrdkpTjZmPs4xGsIdnGw
Jw3ArFDM/U40XmbM77T3imydoSnQfCrStDu28bv3BUfg7Lz2JsIvTdC1/4Mdf0c+MJ+1Iypg4VOy
bvzoB9e5sgnUzo8F52XxXq2aGTDEVU98ErWW1POWADQs6niYoAGjCi9ySxblLu8RUIUtsBEJTfV2
Y4gKUQ4gFWLsCqkCP6HppVPRMTpmft/kL5K/LFZIV1TPKrVlgt1UxPdeFTXXKCg908fzgBQFDqPo
tCvcKKNzl7IEXJvk9BlVo6JeNezGXqdh1S1O4tdiucRa5RRvS+E7x+GJB77PcJV7pBdRKovR0Ftt
3GQ7O5qwRqPAPwo6k/Qw/gSHwg3GsUKinNbQgRiPuTGyWS1gJduVgD/L3DZ7gVkPNxFvka6JUtFR
KH60+5Wv/SMxTspHHz+Arzwz7ZZCPhtfQn/JAD0Ic1mVCrh4JOv2Bs2jmT0/mIVSfOFFmO6cg3j9
qRGjt7XQ0q6LBYtyvB7WebpliF46QNMb5mfHmw+uoCXEKhkSmjLuBiFXxoTgpgdMISBHlbW3DRlX
Q5N9JBBHrWCbeu55gpAt7NyM9EQ6tmAX2cZBu4LduasP+coQVBd3ZdkbLXPFsKciZUoqUdfyoy62
ooICb1oXCrxh0ekI0dW6LEzLtat9c0vGyHUPsNQ+clGudk3oEKFgo8dazaFMgI4XST6+Pb4WbUBo
T9hrzY65MTRXshd9FbBJ1sjbk+6Z8T0FBSZI0fC4rZ3SSfldc79badgs6cSHMPbSTbPDXnWUpndt
kM1GfFIcjJyKU8ukdKRVtyizi5M2ILD1HKumcq79VI1FvkvvMxcuSUPlOeRobPeh8ritYMrjGEAC
46qC9Lp8dqPjqyneW5VG3pd7e8LKp+MycIczWjnOr2AvipJ6jlT5Fi2WwC0lqmLLNCZ0LGR+kyqK
mmOWOdXlWZe3Z7slnHVFq+3qN0+bMFbrXzkc/pjfw04uSjO0VQ7WLK/bkkMDjAjbQyTFFGOK6RH2
OtL+4A4OntZc1zQV9uExlDBjwcP+J/hIQc7pOKp1WEaQIU6E+fu/snElNWlwyPE4cYm0JKCqr//2
kDxmNwnHVHHrbNEwfLX3cQwEAXgrCTakaylMsUa93rzN/UVnLSPbNDYuZFitDczK5UdHFs47fGcG
luI26P+3ayWv3pl6/ZBg65XBKgHqRNuglkMV/lzXuyhWFKhUdW3x7b4hwBZbM9zSq/GTt+WjVny0
MYGSAI+fLsTMH4WlMfTzP/jawXD6TJliy5sFoxz09X3+XXP52pQ8MUkzEZhixoywJ3IXVdBCdqVX
z+1np2LhMxtxkNK4lQIUrjv20lKmQKi+mgEUU1EvW2o7ScKp8CIrFjsVFApoC5eQ5R/LRFU6t1qN
EQ/aLRaXOf/QcWb73wSvz6tsHXN0NdyneubFAn9weCWNyx1Q7InpVwFYl1wHl+Xj5k/d6SlcXi9L
42Z0+JWTp6W5ptcvHhT8jUq9sQrGMHSlVqNbFCl1AXzhl3ci4dRdZLqW8L8/NVSgnQ/wHVisME38
KXTN3DtG5c2bZdLOAWG0UOhHpV49tNk7uzCT4yfEppy1AnuiNiSq+NX1EsV3rLu0QaNVoauDlt6e
owlDVT7CY980c3GonKS5cQ8ZJSYYctyPVc5oD88KYcQrmBxW5tKFcORv9t3NgMrcDhfp7GCxsuE0
TYMGXqtSJ+cwmuOgiemZFhYoGuUZPLP603lJxPvVyM++bIsTY3gTpEmi81seMSOYAhzV+VKQnEw4
BbjeMZ+6Mt1ZxAomVuiPe2R5l6BpRme1aGT5crwBmaz0OG0stZWRkoElEsJ8gH/wyXCP+wJHf0EC
+EoWFbqwIlmrb8YarhaidEqMuEd3FMDvmuqxC3XzXJe9tiwfjIJkyNTBHbEylwrPSNZJIECNRzkd
RnLMLWQ9xI2j3eZPdunYC9ns41oGFAlGBKqZsZQeU0yded6/h+Qu/VfMH94cL/afuuudv0G1VG93
UDPpQ18+BedQkKpcdv+Apimc63MneI88EmfgsrumHAmUCslp21432LdZPo2E2RydJanRgNE3lL1X
dE1snINVj/amdkzf7mn7LGe+cgWTKSdGhPvbhJuHMeyb51Ti83JZdKJt4RXr1d4gDF25f7n2BNEY
KHYunvb3MjHczeksL5gteUhAYlMMysNOiKkPn6PARBWWCOMvdR++ndD7LaoIk7aIfn7GiXWrjwNN
VhH1hYmdtLZ7KqrxJ77iuV9WiuIu4mHT3nuZXVOPU0N+QYrCoWfPQcLZ5yUI3RDUIJM+C72I3w3d
e4o6ZuiE0Gd0iWjZSM9BnQOUf/adJyHvd2Nmz7CYfTRPGHRncqUtRe6Qy5BYY4FmbTCiy7WYvhVj
ezOLCVGaE9cCAB6zVFmHlIPLxHnGarkNeao8hoNW/1azJrLQuDXs7Rgcnzjpow+TBExBSO9Nm0fL
pZuDID+Xs39DzkkJerRp/qNenF/3iULjIhsYOb8KGMc31TChBmXg04W1UL0K2IVV8P6l99UYIs9Y
d3j+mwe8IMq3x9F8ee/ZhhIt7/IM0QEZ57etMSaZOJZC448Cchv2wnmLqgwjR7qxBD3P8yzKPTj/
20hCXTDDTafmUKezSe2xyJH+AGPU8AnzkzfxFGsmUtAp8s+KWhZ7BdqMWqjQrfg9KtH+X3hbY6N/
Daly+NY4zF4lQjc7VuNiYxA0R/vaTAsE5ci6NfbAoEY01rVylFufV9Bt4PoMSkP1uSP62mmKgPvx
1dx7pa0N8FLJM3+4bQQR32Q4Fwi9ieve4Zjfme7+FGFZZVpQ9gscbGeMyet3DELURNQhF4H8YPrv
16QfxyQm/I0ZWb2pOwbWwjBBl6NqaRlOH6CUacG+vMhFslx0DMSM+D4cMTqRnn3rcWnHkjCS3iHz
+juU4GVy1WhF72fjRG8po+vxHc4r5AQgx5EwMxOH2SQmOlWb1CIS3GRyGQSTdhXQQDxDOZ99r6tq
4nhZSTorgSS+bBhfMRJmgfVfc7OmI2TbThLcT+BmLQff/IBvrlNpWmAegtFcKpugbhbs9rIKcX3U
inBKfdG17s0QmlC68yklOawOv8WlFJ496bTRtvAVo/5CvgJ96n8axI8ZonM3DIaB/N+PvWG1fr4j
/5zlXzXYoEVt+WCRhD2oKc5oAZLzHx4TR86ZGqZ83apT1iTUp3uqDZ1onUvcXk6W3UizKW6kmeQm
64DDzXDatvpFyCEb1eUrZ03+/h7Bn69k9PsxfL2mS3dgDlhr7zT9LWyKhdikJs8Fdbyfx4zW2HWj
kzEuP9FYWaZB02RkGxIWQn6XodSXZ1K/N/P+Y7qmThgARfiFb2mFf9LDjl8VyL8ErpEAyiHPDaV/
ZOYH47jhvb8CJGaIu6Qr9JDLTlTcM1twA+hdwexRXS+8UHi08ic2EAdHVOclBpEl6z+3YD5L5HIO
TY7swzBaeI8rGh3JNi1ctBsHcKW+pxejFhzEUSKPvjW23iwhQKeWoy3Vz1mQDW11qDmgS7QDcRu7
LBJetFuPd+KX3DGckmNvzH21yl+ELROV62ngK5DyNqtTQR43Ra2ezRZEfwe8vTfyDDQmOYXY8IrK
jCdlRE3XPeYKmoIofWUeHATWP/1zvYiDN3t1mJKbnzxBvJLSNZXuHBvduzM4NIo5I30q/L4eWXBR
GBArqNUuF+mey2KWsA27ql3plyFIIfLVD/Awekrm0rVVe9pNETSqlPzXri5x/7SdNzEL1d7nMMsz
IzFrODt7phGA3fef5xJysIOOXkEhoAP67aWdaSp/zMnF163EFKoMeHUFRqFml6k6E46oQpnovn4m
YZBp7SwbhSG7S8SzY7q9L6Wqqmf0o1u+hpTfOUBakWDNn/IzMzdOPBngj7jEqT3iemkkeNc5Pe4d
5M2N1NY3ryRbxSaHSO3jxoS2pnaAbJWm4JbMJJHPgcHwNlkT9mICxQyXwssjZkCSaOIOKnEFCwra
d5WX6mTLwDlclDaVB24j1t6Nk3G84Ore1grDTLG7HBqoGlP17+2a1uZ0fKhBcFuvcXnDCIC9pWQh
GpJn5wN1wFh/3osMXV5JykruZA+Zb4rB1LqHk1vGNuv3Xxr8i644AMlTBk3i0YFAFszsR5W3f6fn
WEPO8vVvfTwUOmmotI8/bqUa/ImCrR8usDMCSq7xcMr9+SbdVIzfb84TzMWb+r5q5MJWdHN6oqUN
X6C145/E/C7FCMmqdKRt8xrtsdQ153ot7Rg0f0lIBVUtStrCCHP+9T66tHoxsowhOQihBbRonAlg
tHxoR8Ktdzm9ZJASnawU3OEBDALwSX7MCQfmfvp7zrJWczyg6VdbBlr0EFX5UJyoIpQljkxQtsjy
XPZ/LqPaNNSwYQi+RM5pkglWOwEtgrONGnugXuEOznrtsVMWSLiT3STFpCwhSryL3Ht9QQsiCH/I
2u7rIpSfVroaMqjqhfBL9BV4MdlFM2OQalEFUwgqWW9yvq78ypNYIA7Ww/C0i7fL0d3sV9HrMixM
BKx+eVHYtFFghoRx+qjtpkU6/wouPWEC03aWvJG6LxVv9lUVdQjnGXAF/OUhwNUzhuBPDQIUfKxk
9Aj/klIXwiXjnq3p70a2wDsJgNKAPfFLrrsSVX2dmXE4MzHwKhQFvP25MZXo6+R09/TtMEf/LBs+
SGW6m1PJpHd3yrtE43ba4mgJMZk+kk9M+zthEiGNV+fGrhEa6EZWuYa47TVu4ztwjsjj+lM3yFTC
QdMIJV06tN7zwNSW46EJEOw8PkQRjld2myEFhwXId1qqFgJfsaVVn7efW0uM46iy3C6Ph2E/Uq0D
MUAP6Ht2/+WlhEis3HNYuofuzDX7vctNrjgVOY/U+jvlfmajnBwv+fbqgon97+BVSH2+5yqBtCvY
Z9TSxrqEC2y1eBG6j1caUx/AEHyQlckkrRvLc+2YDRtziW3+ABBAVCbwT0zW86bS9X8KZ/EE2Fxh
K5rdbfKcKQyFln+Uym9j0S3n55O4ATcScPUH6u26kG5wUur52ENvPWvUbVODNMVOTatiC/9wk9u0
dZHDi8B0u5nERG4ijKK7xL9C++YNBuHDFPdy5I9jig7V474crzB3B1Z0GSlzYdaWb0FS51qj287N
ASWwBymyf/tOBr/+Q8eUBqwo4L98cDqTvOUQ8qrThlstpId9BiHaWaGU/5WAzkwblB1H80bE2yr/
lRWKygA+fmpAix5cRfCHa/xZzkXBSfWPHi7tsUfWrcDsUIiZuf+MngzmLw96It25eRmVH2m7GKoQ
zR+ia3YI96+MXg78zE0xAPi/ym73ONd8+wOIuxSPc4gzTXCTXgYmVCw4+HjZPG2qgfZ4UmbKBh6v
KJykG2sWeDCJqDLDKc/+Ql5wUFannB2COAAkHJlSpkubgDh8+28JoOxBkNozeMoHoHwozBnidP5K
vemaPgCuyQEX81W1xWJe6qJinLrjKzV/Fxo+C9GNbe5MUqNadw23zV87eMS4UkywiHV1hW4t8Lb3
+vJPTCARnNuS/497lxibd380LqqmQoZBAezQYTs94wA3xkdyaqHMhS4sSgl1H8oWRiEvOeH6fWGR
dTA6MZ/7+QSiS2LuFV+RVNi2ggi07XXYHUYb0v9eWkCoDemTSmevnslcsPHKRGcShZANCcuHV1aT
38ZrZS0HfTK3k2x5Lq/Avi/fD/iZOh8MpWZEifJZaaH1ZsSroPUhbJ3FdqCwRPB30xcsLZBOQD1k
ojMAT0WVk2yrwDjf0N3Ywikekk5T59rKqf3F9t3qoUfugTL46Zbv0xHVQ2mkUNCehMhoBtsveFCQ
C2KDchZY5xUXxmJGJOcCCoVKXIcXpGgmcftBHpETsSOt1VaNLB8+nbQNj66RylbxAfFsBcdPSk+O
7vBusNHAs9WciIXWN8WyJHSej5eB3PNlEyBfLRHxDFPHRRVRUWFitAsT1C2hrmFuU9oyVUo0VuMQ
29uxpd8Ecrcv9FUV/zb0LXz4YqtT+mUvUfZG7IHDJdITmIpoEAn8aqaLy2YTQM/uHq5ZeDO1QgHs
m+/IdiEC2pdmZBz9nsr/dKZ8JfKW/0j+bo5XJwTibjdEejaC48QA9vZgT/OMrdyq/9eCUihW4IkE
fyP9rlxuq3tCgIpYozh/5smuTsG5KxIJQ3w5t+einYsCDdBhxgT200pzHiF+TKzr2s+croaz61zH
rokouR9xQ/QPkRZ7XN+m/uqVFL3z1Cx0Ufg/n2bvwzjEff0rCOGwCyXihTBsnOwDHmZMmxTkKoZJ
HVUu6YyXt53wBdejxlebiQ+nLGFIBNf6Yx3E+ArRNK4I05rW1PrjptiItE7gZMtUd5uJViBHFqnb
CCfhywlcn9gWnDlDG+hMuTfyVTThkeDuvW4F6LiJIncB+7OO8c5Ep1yVtmpNN2d3D7oXW5RUPa53
d83RMtztdgRLsD6/Ffn5PcU+aQZtJqEvzklDVDTf/pXfF6eOPjvQSgv7/Z52rpoHmCGqIte8KeZ5
vIq5VUstHVoSFf5xVcnZpJphf+H8aVuYGy4xR/IEtSvnG2kPpubHywJoLMsZ5R1CWfdW7pbfOAAN
oke875PElTTlSBWUJOpea4GZP8yytyWF/7mM68jko6sR5kvxQ617I0aT5OGJVlrcGhvAkvFCv54K
LG4/M0HEFAtjsjzoG3Jl/TTTzzEgDNvpd9KEk+2+quS/l4C/qqjc18VWLbgJtUanVKg0NDg+MDMi
sTUtMDrhNkO9Z+smEpmnWxlL4B1IGXw/hA6KwYB1c3x3tkZOM7zfKYlcj2w2R6o5bz3vj4guI0oP
tfJgZ/tHI3jBYLJ4IUXvukhqdjRbVpYkk4o/b301eQxDYUMJfiucJT8IZ8cO4VC/PqiyUFDYlZ+m
NPuBzIOE8QFYuigaf/5gYP68xoYqKZKtfCc31+9wlq5ca14YcdZG8J/cnG5/osmChXBfp6IyM3d0
AdRmHi55/LtAPhuaepyZ8y3alLhS1hWpriOZ82VKjVB2UlcD2wKjcbHnXbGFHHtQ2AGpC6zdQkPe
dA5u5Lg8TyHForp/RlVA5unhdeLU/hcd7GsfwZJ50XPWDI2zn70ELguVnY6OR2mx7fcWEwVLT1p6
JB41rHPMk/9yoQIMo3Ngepe59133CDwBgKs/u0BL3ghMsgtawxX/2aAim/I/e+Eaydx/YSPyAd+s
fzHSHJJrbda3DVCGCYVg7nysxwgB0YSIHjcKxUcpB4FWX/C63Pti4mj1jdIX6PXTuPNKq7igbFQC
37bom3d4b3M0oD2SFpz9bY0y1n50b6n7wgGTmA9vbOmh/UApsBIdSPS8KlsuHvN4COYI3+b2caRT
vmh2m/L41yrOmdSfU0GE+2KVEMfMD9W0v71sJc2szMHp9bgtKd357BEIGFgKkOHD/QEX9NDGri0a
Wwjke12Wr052Gv2Y53Qw7g8p2jfGVR6BobBuNkYVhR7EIf8iw3iO2miLmRpzrwGJTM5w17DPs47I
EJlkeq+W8Vw+3b2WeFCCoi3sVSLAU/3ZhP1y4E0DurtoL/JFHBc0TuUDZC3gRku3D0lWXAiGpORh
FuDd2xCi+Z2z49GJYEelw39HNeJjEMlE9UsLE8f7neK/jpombm6p6CJzsvhAh9yc6XE3A+BPnFeG
X5xqRuNBj2C4JgyMojdzsHluSTKALbbRTgmv56urpoUsBFZQfwJvQyVKptL++B9HXfodvlLvjmna
EihmdtBfYoqTLbuBN4jdpYrDbUr7RPbM7AiWeWjzRtV3SQflXPIKKsDjirUV9apCdUiX6OQvk0rP
gvQBmmvyhWl5b6pZm0tz9xAQl7WIgf1Odg2hHsSUDqMeOOHXLMpcflpvziwEecspX+WiFhRvbFHQ
dwpUzu2P+hDOqTVw1vtyKNATMQsiF1j5d/aTXo+fCqv3pwiqFcp3wFMX7QAiDMv68Ss5OC5DX7CF
+wsWAVa2QVSYO80sSYddri3/lbhBPITsk3kd0o1zMNdBLXPtOgLPu/NZ6CQtPmRgLd194cW+J71B
BOdfD1nTZLGKNzBoclITMps5CW/VbriLTx8xXLmDdpK8+M00sK5OF7G5UtVP+pfchW+Lk1Xa5cc/
Mra0BYmRSsS81mIl6vsOWoN3WIyg+ee5BQVWt3WLU/ezixfC73vl6SbK3FOfqx34r91CVbzsr/h+
v2HymHip7cjVuss5pQX8KAKYUjmLpiuKB/5ANhpgbkKI2gCV0xNdtBiONTtgxR+fmpkKJ0bggB51
IZdIjP+OLT+0hSkoosPCMV+IkD6pNHxGMgMdfMeSdVjtTNV4JWGadWizdamdRscwgYhSHNDG2acv
1OjRXGgGYdE6HF+P4z+wpByvooZCW5PKyLgOKV0cygqyJBJkNjDM7HcVHKlovqkEDjnvpkT1ygsQ
anbecFRVwNkA5RJ7EQ8D5zkJgUrRB04bqzK+iKsr8D7t40uC8N8Z/Sjn8xO3efutiRBPsmyf8Hlr
x33nW1EH6D5DzAl/xnaMxVhvefuEMeP1BWMOq86nB/1QdZPhmGj2e3C2o4g8ZOrxH2XVCZ2ryNGn
wlr4LM8mUrmn+yUBZu56dUqxGUCdXK9B0Zm3B2CbqcY7HTm/SPOk36VhEU8JxP2Bq703l+VbFP/+
mbbrSu9Y5CS//6Pxs27Kz6pS+E6n6n6h975vFN7zbbAnBtgdWHu62dLtUsepCFcti3igpB3ziOM+
i1jdHjmZ4Q1NZe9CwWnSBhlosGfJgRZRamiE02MzdTF6KXzSgdDVSU6gTyCHFquHn2/M7Yu2sVMB
BzME4Lk/W+rnsxe4c10y0LSNYvOcMfybIUR+NTvyVSXYWehUty60k9o9fuLrMkhzq4EjwxDh99Js
v/HWLLlm2C+PnvCmHBdWW3Gp6RWkXeg92ZatThv24cLE1GiC2EyySK1g6bclgDvvk0Tl5boC2M60
cMT+kV19AHK8tghjR7qZmNyiZdsMOVZIBSp0bk9E9wbS2U3C88MVLRvZ3KQFfKAts1z2MxTbNbv4
bqDYkzXW6Ucfh+UzE+XcRv4MmAy1bRjwn6iz2gRsThz9E/hECvCkyi0FpmGAMffWbOGByPUMjBud
XhNcsKQkCnozyANJmMvxW7+Gu7HFfScfcTn5C2WV+583VqyIUEJ2UnXz/zDp2jqN8rhPM8pLeUAt
eWh+HtH9B5+QLqJS+0I97X4WmAoIzou1e3cKBHU05VCfzsdOeF0dNWef92IEARMR0zrg8Yiyk2xQ
11pLBNJg1ZmBVxi1SNJiczfj9/Wp2pWGKcCwo6tlZvwjT/ApFeq5Ej3ZGRl4L9oU4KoaiSoK/6FD
usKuGDBMum3j9T0NclP0SqMoNEcvtiFBg5G0S52vD29gNjX2omHc9bEW7/yH/3ba2z9/Qmzhh1N1
P6ROyDWPjembHEOe0Uk+DsFpjW/Wg7B+p+ERCZ1cCEXvRafc5wd+Z56XdZuJZbYsteRTJ5VtqD91
5KdsPhb5e5Vh8uK6I2jWf3Yekk/7tCGEndnANGCLMx152pwdr9Do/J26/cKX+SGxROreOhR/pn9A
zUGL9W/RFiu/Jxd3xtPO6xE/Ow5FrwgeaXSRtG5QtWegB9ElEoF6oGN3l/Frd4ufHakiYKQCns7n
crY5h/XB6YPLyl4Q+7JHPL3PRVV+/A7tCDb5nv93oMAilC0OeqUfvQOGh6QwPvy1vR7sRcmid1GF
NVZ9V6sa1zyqRXPRwGh27Nco8j+3fljQbaf3FFEXsAoDzUnlSUil8mLxckeqO/0mPQkgARJ/hFvn
M2op7p81SxdQJi2iTQGPGNbnm24qhEZjJ2yh6LFQfirylTq0EcSMA2z5/MNwPZgJ5YA1TvLdR+NJ
KIQNjcZKO2kc+b3nvA8tfzPNWeA71AKkKlOYF5WGtOGABAGmLmTZiDqGG8QsJhT9v85R6WscXhvL
S/qF+I6dbGAuXLDC7mwBSguc8/NhWQ8gPRcd8mM14HK4vgE9oDR/Qf0Ek6lao6vQMsrulJD7r4v0
YihdIoNUTnPo+rRdNHVqG5wbe4sovr3Dkg1G7cehjugQBJW9jSUGop6x2QumuSBDpTRxIE6ysk9H
DFC0bgP3Jfc3bPIX+eFv0/XCD+9HmvRwEnAQfuME4e62bgfU0QxTo90TwzX+zivhocABH/tqyw9b
QSBPnF9csO0/3oGUxfngOWv3L0qJBjpA159I93N059C8CQC/d1p6yHwd5PtVpf0i/6DwPlu8Hhm4
XNSYTY+kzf+Ko84mdUhkx43/0+EMOC0neqQtaFuE52ucLOaobwJtCOjnBG8YKLuQ9ogRnLvMsclq
LgeJ/0cxHe11jSD9hfgZ+eAprO1cUkdg0hl9P9hd/LT9V3TmjdlHMvEtUnPxIvXn8OQ2d9mw1Yf2
kT8JBlSSkFnDOQwi3xfMRrUwfvbL/R3tWmZLtnYH1hvfhrVpmW8CzxgdB9bgoWQuDzWk7JvbdKql
71lEi9fbGzLY9KIxn40t6BfZ13msP3DG8im14ZRjpMyp20SCwMnKKTp3g9YXkLe2lp1aAjhII/QH
zwm0QE25me0E04IrtWmmJ6lTuModnXWheE1+Tk4R981JfmF12YCrFo3uyHer2i078Eacc3Hd6lLa
bfQNnZyJcQkXJazFzJkNpdKtPtBwDp9NNsDGVQ4Ky7kn3M80/5DEyqhhtE8xYOoaZABDytDrARdl
0BgTMgCGUhBUHLY5aBOxuSvNlQEanM6drKsRDxKs9afTmjEHUWdfM2gYxszlbLqiZROaF+ihZvIf
f51G1XBMZCpo+q/0ccE8QYvS8d3n0TubKeObCdX6rSBEEfNagw6zj0RAyuh7IjIvjRUdpvbCVUY4
wXfRg76wI1HHvBjftFQLrXGMdjotte9QujREe2WPc9o5gBElTcf3QYYo26KnUNmwBgbDCjW+k8rj
XViSXMaAsLZliPe7581dBfVGFdK3LxAV0OrX8eEjawhWPNw67LGDhyrrAOp1dClQ0mfZfAhcwn7l
QIK3y0t1mwOzmmLV3dKGp37hSx+vGhtQdVR0V0pr50PKGb9aObmGRv3YIL7Z2wOVCGX+8uK67I9Q
HFud9c3oJ0g/IWf6SJe432JI9fr2ZdLhnUVu0HoiVQn8btgSYjlLMPG3LBC0mKAiDleoFxfYxn4N
UJWHY9qHYZU6jYlFNVBNJqB9H4FaUtbPeM+vvy7Nh5H7C3DcKZdWfwHDAuIu5Zd6Y0m1PI/f3Ukt
7y9H2ldodjk42oIcVFpm8Jn3k7lGQBo2d/bO+M0P4VTYFs4dEDNW8vVEG9X98ghymS2+r3MbdFWW
PVXC3BMUxKS9XPjTV86zbUXq4LLRi/l/5lVLyx4UzNU5cvYvub4E3JDnthZDh6HvBJAUxy8/3MNS
t8BnvQVAzWOlEjCq58doJbCWAscULeU9SSwiaK0vqxJykolTjrMdSYNGWImV7iwVVzuXNRsxYDaf
6jIbJ+JvPvWvWEefKpg6VS3kxni/lBj9rTfUoaZ+UWbWw7bTTn/qok1A70cp1TGo0vSaKhiBSrQm
fg8xSITjFzGJIZbqDbNSOEcaEdxdEvmxZ51Po4K/7NdhMy9RqUUiwMam/+xiKWhScOoIyy7jEx+Q
BSgRCZMXq6oIp3SwM6o5Al5fstIDFTGP5eP0/SRT0CHWVWxybaKgz7U1b3QlYXAPgmDNHXxW0mXy
+LyIR9kN+9wgC/EGNKkggYqyyA4aU+kzGM1TDOGlzmXuvgq4cLdx2zA708vFGF7WyiSrHS/ho1h/
eIfDeUWvg2z+/GbqyfzFm/d4gXndAbtu7FnbAeu4sVZAX89Nf9oB0QyCQHAOz/0ERwb1alnzjEwj
dp7aQejs/ixWrs5IyPKMgZ2d7JAwpYJw4/MV3SLuoHOA17OOWBl+ZWyPgEwy9PawTcfv9vRWEOxp
CQe2ZIYpBY/LDPxeFu2kic7IT5BtN5eXB2xcJBD3ugLlB0/Bg7R55sOuvbNulYjjsG9j+7i3o44O
wRIA7w8v8v8I55dmK0AYriS1zjpfARMEDMA5nKle6LvGbBi7EXHkIFyaskrTSHsDst9iGXlnn4Iq
iPUFBaBdOTMJoU1kqIuj/vOZRRR1CuxsE+VRVyZuMFqTqKTVKyx7MzTAcAuLT/97SeDV3JIPJusY
jgyDVk1D4zm94HH2npi6WVOloUCtj/zpYv2sCd6e4AH0wbrqQZgA3reePxlfFvjD9jF+HtoJimBy
5AFgReg3eD0nFRkodzvTwV35UOt1vUmiVLpv8W/k007vl6hbl04bbET/D4jJqYakIn6/X9AWhbSy
z7cxSWAH9Wv00VWT7gc9MYJ/Z5sObSePQsXaVIWvAjo8aAkBlt0I4IQkhOvEIOUa25pZcJSw7vSw
oY96ZrIV+Mo/twcXqCYUW0FF8b719VdDIGjaACkl8njiSFVsJPie01nACR/PVtfOiGLucNeAEnmA
4cY8Rmt/4Vpb5yYdDs5GprLnfF6j1RmGo2SNk0e7pSa3RqfcOYCX2ZR5exnzKHoum65oDZ7YkZz2
XtaFtppUr5y28+GH2xBF4MN6xm4uORuOT+7v4lSLkDUWuv8ycf91o6cYdESSzRKOoBYhe7IEmXsr
Kq7Rxh3hmdCkNDGtJ4INhQ4ukBVrlf1lDZc2p32mrzRUO2vwVehM62IalkWeaSeFj9yjRAnx0I7S
CcTLSOg7fqNEe2PFM05IMi0iCHUtaE5FYtQsgmOXLy6AYJHr35IF4LTC7BlUUSq/+0HmombovDCI
5mrnqnZJV2TwKe3aIlpSV/eJoyYuGYphXv9ua1Ci1eJ86VAnTkqNX/XPzfnADE8iALQYvtBnL8N0
rhsYK8e2zR1WJ6bFfDlp6V1DfqGMJHemlMbgmjAejUA+8trH//xRafvjHRLs87ib4vC4UQTZp4gP
6gNeC56NvT8STly3J5ROcrJuP5Y0ic4lCC09flF283kS/umu93acn7g8Ttjuzk6JzDZAVt7TWwkB
xC6jVlVZlvn/bJn5aVB38T02VJdv5HFs6fwjhS7lmeYP/OVfPp7tCAePB8Sh2qAB0LsgUN+a2M+m
ENLBM3LpAhhJTcJGGgUDsIcivUGCbliGBykM2+W+MRZff4QUhh29VNq+IEJ/J+zZuRqxnMsXfdgM
rIsQ2jyjEcVifiXLeTDcRh8yCv3ZgbKH9fXO4MMMlQgrx9UVE9W/u7vxs7uISb0Hm3g4PVahvX8R
b90WV3gztjIV3hYFOOU56EIF2RZuwMzWY2218mf+OyA/pchldiQPyaPWPGC9cIbioIzjs4kGSG6w
fssIyAqnwWwbdhTd2qjQ7Y4o0nGweKydD9tsSIK4H8Ro8wnaOsFnNskMRBOu0BVr8un0G/faAC5K
d64b8CS2moJyK63r5YgBoZY1eMm3XklvPib8TbTc0ZVXdn+mKECCY59hF9vmAY2M8gioPf+Vtrng
OIqtxBIRE3CK5IiehRAXGlqt4XIHP9ihBGUZBvBtkj/fYNO17Zkw4eNmBDknwhNEmEcvYNcko3Id
oAY6sDhqDuqHhioqrfwANvk2h3q822vWXsabBaW+y9QMp+Aam2E3hf6ICPGD5aDmyRzvL6kEqbUm
588G73oWmzxNuUKGvkpTUsIlyJDjpfeO/n8LpqklPrJ8bOXWXLq+HLz4EHZAIIKuITz3ZI+KquDH
+5oMVh9cSdhh1TUFOv9+UdLXq+8ObErub/FbXdLTg1nfUgAuAiwSYTGIJZYeyffaLnPjetBwZ8Vx
pkrWyL1owX+yVgN1k9iHpL4MUQpKnu9Ltjwodd4F9GsQvZ7GXK+QTlo3QCl9NnVBOv7eA3ysEOOA
h0lfbPh11y7sHFWyrjDlKR6Ob9pspQUdJSjwgLRTmYTFIgtaW4aObCiOcyQM9YbaSlxASCQJAQCq
KyEjTdlFpMsZhRq1zgsXNWcSbsBlLxUdbsUQLces3COeBD+mgxN7cDkCqJP6SDscmLJzauD52bfV
E5GZzI+ZY4dy406LMaQWQxOO+JPkFHiVFdj2n4jJhjj9GgERndayUkBSEP0B5xgkDnolYLkp4nQY
HHl27URS8MLvHUCM0t9VmbHFZdyPgVuF1zHWIRJljyLeANOK4L0eI9yOieQ3wOjapcbbReTWUe6G
EYr3iYEft9/BYILUv9cuh39y1QJtFm0wJ9+j2CrpHf4vIonEXeIvM+mLHzuCrSzJjvt0OY0zjldL
B0aO3C6x3YbqF90CC+8CwjSPU+PQ16iez9hJyQuZGat3saHx+/XbeQHA7JdF7orh1hvO8x8rkVS3
9M+ADVvmY0DpW1cRKRdpB7rn+d5pe4oxY6VxfcTlOLPAhUO7+gNOLNJ94hQxDmbzoJDVQR3p41VG
tCozZ3NjRKY9JU2EwULiAGlQdV23dc4ddFTPdc68PCJmfYXGw8MOamvnr4uD7h7fe841I+hRx9m6
F8HhdE17UctyWWbC6mC5XXUENw9J2trFsunfUtt5XJ1JQyHGvzpWTwkwBGChnUSRKLbZDRvGW0wf
cHFaiFcFJvTRtJ030VcAq7gaQNT3qMYa2Ldj/9MLpRWai3hNg4euJZQkChQ/ayoyb9wJbQy0bOK9
vhGOndlCsE4FRwUVE6y+qAnMsmQQL/bn/foTvE1Z7m+rvIqco8u6ZwQ1FA9ddwXace1HOVPXWjmg
5l4hemoTVrRAfYQ306hw/ihDNAx3szcebrWr+Uc5iZE4Cz4yVIsM7EcAQiKGMuquESDD6jGSkUGn
xruHUNhWqZmcuQn7+pOBbUikTThXfRYCkfe4bbsf4eljP3WIr336z18pjU3yCuC+q7CC588KX46K
e+i1Pq8crGQPOwqcC8j83FSQJJ3RnrJvX2ElyvDQZDeuXSfW0zcKaVwDYT8kNMVd1P4G2kvk+hvA
vb5hxLAvmj3xYfyK+CxyUjlj7B/n0C/zkqEdhV2MvkB+ab0+XSVI161AT/2qMetYmrQ5P1JPQdpF
+PTG6kOT6QKF77jScQRlp/3U0m64MSsPADpb08u2avdlWo+k/YGHMLFY6i2OgKwVoDnQPg5XaSQY
YwO3+xLQYvrJ+6WjG8p0/yRk/LcVz0IlqC62XUmnm29JBH5x6nELQDKTR+wt+U2d5Nqvf0DvoLza
8JA/ODJih9QlvspMkOtK493ulVwFRUo4QIaB7/HnOloIDivb4np6T+ew4mUtTSNogQVzSSyBNw+X
hVh161su9Oj9HEoBuK/Wb/YGP5xIqaB7c5u6KzhisuqBEgqXNjSOBsa3b8NMqimIwx9hw2GB/bsD
ZNv+ClrKdKAta/7ht+iqF9DxVV8pjMtDWieL1b1F9NqEBC96CjfRaCwzzH4umxjEu3374ow7oFzO
fIYoiy8LQ9TVs06evgFW6R5ix4Ia+GMFxtm45t3VRXJaoG5GHmwep7+Za+Xw/oNPLgxwyQqClz78
Cj+GgUrjNPLO2QBaopTBviV1aD01rCNWaXaLCOLoG0vKrNV7Tv/mtKrNkLoaCOShlNotZqIarIW6
X185cpb4tN6OHIbSTlKU8FfMq9K3Uu8Kqg2rMP+LZkmYSeofbUFaXV7rdVr2QXVJ6vIGsaVl/Sr/
X4ZJJdPRgEeP5bG9EUSs/42mVfoFGBllQxIqoxG607UAc4HZlkjOl9soB9WHZaJ7j46D71/Xy3gf
7tO0L9EGnQ9efLQ0DQRsBWw9+veHYLZvFrh17Eely0QHdEviBdjDU7eM+iKTqZvL3DGtsDY9Tr2t
E7dW1uBlvc7d3VaCbetX90dk+wm+N2R43KaGIUq9RcOy0b+bBa7XEiDavIwjikjoPSqDG1JQsTts
6Bi4KOJrTjfJ899lB06GWx4kZSY0oieUxywQwneTw4jP7XDhApVJhruw1NuI18d4uRmpiAq4q6SU
lwZCFoDGfvHH2VsAbG8nOZ7lOcw+/V4q0kRC50bhh7iZ39yakTq1kHAm6+nRedRTEL9Y+PILtORh
1IAhLyzPpA1JkwYeVRxIK7Y8bFoKeo9yU4DZrZ4YPRBmtGLJ8Kh3DBEI1LOFyzmEonxarfrEXWqx
YTCP9C2cFtd+upWEIIH1V6AIWByI2OQlMOJKWAbdy9DNjmZSnX85Fc1oGQWvZd+kCsyJ9EMV1yDU
lmOhKJauzr/dHsZxjT78UHd+TxLWC42Uu4znkHgPPcy08TtONsMxzCqxIBRSSuvwCdzNzWv04pNJ
PB/A3Vl9G3dJ4iT6VXffMEYPz7kbBR6W2NxeWFiWHN9xVjepG1TLjGQCZNTEGBpve7RGnjAYVmKE
oKVeFJ51ATJ0hxcackV9H7/c/fAQh/axuOqZkrySAiyFe3BTWvzMPmhg3eC/KmvqCV8GSDtFgo+P
MBw237FhyVLBHkU5Np09uX/eOQ5dhB92wIcHcimmMEcyqduiiVFTVuslpcp3pqZGXJJUdEQkj4yz
gFXmBv8/qyr4aK5rRxX5xr8cTVgH9A/GvzBJLYgoA3DV5L3oc9sr1Tbf/4bbH1U/pq3VW0+vA/Og
rsvJl6N5m3Z/OZkstZ90sB5mERQDN8tykj3lmYXJ+hHSfzlTR0ZvPdb2jNm0w7EGbfuJduP6+34s
jFKNvihFVYnWJ+wlFgvysJxm4R1WjX4LyE9BJdMH4YFukhscWyGX7TsMILSrL/Vg9gbnbwg/Gow2
NZOf/28fXhu7bsvn1BWUkoiuWFHPbmeY842O7Qsy8YSyWr7gdQZRAyPjAehSRjHWvoQCZC5Nuv5d
nLO4nfqoviKkjLaxzWgyXUmeQBUzIbfKXnTJtAw+XA1r51SLHhEPvTauAo/Lbocp3g5d27eBRCFi
Ned1laV47m8QhgEeHW8uQC+qPH1ixIVpdYzKk+R9XkrOQdIo53cdxO+fWED9tyZ9/YP+yDKIuaUz
FZZ6WTvTPEidlNN6zjDcjN0MJHx+kPIQC+khnwVndOMTIt/Kol68fmmendf0ksia05H13SOSOgQF
frBliO1lDnaXup4UtSckED5NHRGA0IQTgEbB/bgHG5cITNyH1Hx0W4mGnUKvY3lLN2kMm4Gf96a/
fXk8cYTPUbTla4IGjKnUqJwAiEFqX4FfP0+g7nFow2YA84FwTHWwaEpXk45dKlMrxmhEiyWgPx1E
7XvVGpfnpqWnXBh8tnsVWEg1TxrmaqPOF9ORbMzPn3pPqNdcQtSB/h4vecKcjKQZL9CNRhOa9G7a
oYJl/4LaoBsuKfhKD+nhthXtzEqVHrrqqWprCcOqXo0kc4cChbJgIqdbC8iF5t/n1br9gV/q4NxI
udCoTFpQB17x490qDgmNXbbELLiU/UddzkE5nB2H6Hs8vNOZmViOZB8XzHTPeestS8cTlFOTbzNN
IjqoWVHLZi1sPhiY7uop8pos+5oVhquATTCnX1zo6Ln7kE1z/y6SYUR895qDe/sR1dcqcSpjZqDo
tP5hF3lqJHjv/+Z6Je+L93AEVsRTn38NHSa8tzmr9s/uQXAExs13wQeuBHmjvBnniYBTRJhtF2mx
jkzwfI2l1enj/BsndV16DUuvV5fvFYX5OT2c85SqCCYcQLuC08arlUXgEsT2xxZ0tIxFEgbOSFvd
kSgKTRWGaP1rG0A2kjDxqx++bfPvbhiGNkCNWpUV1AjQJzHwf0wQkDlsihO8df35PhH3vMXtfpv3
rwZhD4ulATnUOno/gZBcrd31II62rIvVC0BGG8eQW3Z35eSd4J4mNT1C5tAgqnUfPzb18UfUEWBr
FZ8ikhoiYX/H2sCpNGODwoMSaspnvCHmoLExj9qHqr5otK0kTKjtZRz12JwmEqfVlD0G/KPWNCY9
Uj5RlK4lhJCwmvW3wwAAWnNAA6D+60vvhXL7p+jqryIyDD5gfY/l/T9LO6gVQI1yMG2siJ6bk7dR
sWMlpBWVrDwvRQLeeyb45jWuCmxKZsJx9kzLYe5Vvj4kCxWdgejjyIF7Cr/VLDGp20btpLUwCuA7
xBGE0ONZns7sQrX7KT4nrRWsOpyH93o/J8VpbHFaK6SaEf64IKQwx7I1O/+Isi8GaH7p9dp9EbLm
kfBlgLwwkX3K5negMesDF9MkxWiGoLOnV+m/Ye7ka+1heWtTNrFvNTFd6Ih1XQPtd4X1IHLZ5PhU
qugiSFyI7qd95FjINfKqoHM7vIuH9lm7EspTL1uaUMRms9Osi7EAvAH36wnG5ODgKxiaWftMn1eN
/PJ5Mzkdt8mN1erLYuN7kYu3zUV5+hLj3wdeJi8Rn5IN0QImLO4X4WMknGHkq8lZzVL9oWrC2+2U
jsC5g/4h3fTL0XfdoG0uSbjLJ84EboY5qI3UjXJ73pZcUGrb10cYYQ4x157w1hb70AoqeP8/tyw8
Jau0xNgCYjmDXbOFObacAo1dm2z0u99AXYrixm/Noahwh3R6bglLizHkAqMBEjQ2+h+8kyLLi2tr
FI7Y50tbtKfBjVXE0tHn8tn4KjINeF1YEnQlYewmWuRc7F+ykpoiRrkjzDLFMnClF4C/u92B1Zq6
u0fe2jesyXq2QOjo6qkviHrB4PxkIjrbY/cPGeYA93m1zwZvJZwX5SfMMypskTeFXsh3oaVy8lxN
nHBnc6MkGIrmtTKtbIGSNQFxk0R0kq8qPMLnOUi77sOpnP5BqRiPKIheJDAyUEb6ebJ/lzXmtCRQ
Fqt6vlLTcu7V+f4A+dffNNd8SfDBQBbaDir/gBLsFz7XqqINznYRUCRWQLlDa4ooa+RMaskRv/hI
LEKKPKDqBe4tIdf0YhJT0eTvO5YvJxI8nlZ1crHBkQm+aHqRzU6FY1qfI1aA1Iw6xArM+00kzkIX
BA1Q8gKXJOkgXFEpv/Uv1OdXHTmRogU5Z5FSFLRLLItp4qEbX2GwZDV/3fvU0UxxR78fbBHRGDKC
39a6X3o1/ZGnxu6RpnE/7O8QG2bWqimF2eCuQtd8CQsSHM8Lmcd2XQdvK3sgXSXWzjjuHvU128eA
f3w21Nm3UbzlQ/Zmz5yScUGCHqQMUkqExm/4X3pBLrchP3SnqW8LYIo2Ol0JkIyu5jTY/Fz5gC10
ebmKd4J4Qc4n0MsFlc+NjgPcZXWEI+iUziHdmU4ejJp+w+SQjfvbTOdnNn8uKHF8ZqHUCze0MGDe
N+7Oag2Iw7CRPnLhE/0yS9PzNTX2Nwy6Eu/vs+RNi5mTud8TF9+4jC7AiTJpOdRTUTPhUurKh/j+
N93Xe7sXNi9nMQENyl2pV2A4IIP594G+kiN/P2N66MnQl9fqxI8G0hEHIBBpZLkFr6ML7BzkyDpy
tVuVt0QDT9tkBHM6L9k3BOvnMeuE5F47EDKTbbukbGepUcmDG55NGeMIljD0V1sxJhBhMHzw5xp6
CzxBJYDYgThqMH/UUb0vd8pQ3SWSzHvXKImEr53PcF/aoV8j36TSjwcrTyv9ukZ7EkTpmtgk0mPR
qYcpfCpcngKVBLsIhPLsONmdVLBFAFjeyD0iFS9dQpvNK1ETlz7eB8sQkuFagxfxlVaMOn7tCRSy
RiVDyc9CnYWhfiKD5s04ayTScff537itiT0X4yKkTo40KK0LrpbjDLMane9vcSiR78hg03OS0tWI
9zjpSyuayaP1eWhapZzfgDDF+RtQEpNPnnKAQuQaYcSQSFSiyOnn+ICwP6t71CPjMbr4Ny6Z5Rw7
Wqql3JHNuhxxRw88LXvHBMYoDzmdoIVbqMoUNTSnerdicrMMlGNEahyG7liST/+XB/grLvHTzmPb
aD8gzXO/D1WqBi6maqd28MeyXPsfN4vb+uiV7pZDIyRal8RYlP3ccQ/dVBVi94AGc2lEIAZbIjIO
ChIok6AVg9jTT9HL4bSYbU7ykz2DBq+9VneXkXKx7GnH7fl+KtEN6fXRFMqjXuDqwaAqCyw4l5yo
YGi0+xbm76yIpyUFtZoMIePd+8ipUh3/c7RHDX5AYbJ8cxM5rlRhAHw0PFmAIXF37ZPil9wNKmzW
SNR2nOMb2zwt2zlKHZlKe8D3GtCQf7HCi/KxL6PA9ZrJWjgXL4Q2ni6sydG0JNcr8PLo37tO74cV
QLvK4duU3uJ1Zzfx6OV0Ns7BI58mBhI4kov4RUl4efVFSSF1MUXeWVWuY/Tiw05+07Z+Xz5A40Vr
RL3lgzPbhIVaIIO+0StKsxzFXrt+vVAH1LVa9o/Um9BZzqObRyPKnNr9XBoPsXfaRRuXwbPrVGTH
9CstDFBMkHw53bL1IOefFXE2u42RBQjFyICwqm6VJy1VslmPye8qgBgHRuHhzBhoqIbUflmjKdDm
Tr0TFceWm6oJTi1/V3wJuRNen94hUAqH2W5R2zEi7+jAaYgDkhMzx3uxxXdwcBh1FlDxFc3mNCCy
NnMt0FHpNIU3PwD3IVfROM0V+NU8f0sqQ3P2F3osf3imvzW0lpMs6aVSDpOc/hPM+seMKb6exiIg
HntKjLIip/By7VFh6QLNH+gpL9zGkytv6WcPrScCVxHgrqr6sY/B98Jiu8ZCE9oIcfcBYg8+/r1v
GH3fv8aIlexlMFUap0culdFkKYLAt7VnJIV4mZOV1Zyt1EWUYqqNpKdRyKjwKfbEASBJivgZFN0W
UNU3TJ8UxKVOhLpIWE1L1LemQOjBsf6itSuTHsLtEJYyI09f/ShEOwKtM427R0dI3/wJKK2tSeUF
HPBOgFQzH++khwwiXAAD+m83mkuyDI52h/EzsuqfLgJp5xso9vH0KMDPEx43CWSQJWAER2asC7gG
XJ74+EcYD6EZsKXIhsSgXnZv2oGWTqhLi08pr90EphFJNlf8lanHf6/kPZBnXQXv/IDqROsg2t73
x7t2untpoqkdAPLjuBQxPLUrOYcMqP3Y4ftIHb8CRpfD8qF3ibEyF0/f+SUb9tOOw51KoeTe8qtD
N4upEeBgba/3ivKyzVGrHd73KrwhRVj6jsbX9KRxg+IFApG1uv6eCoTz/V7v09DIFWLz8yS1q/zq
g7Fai4IIqoCVv2tUwABkuHnbAHNfwNt7OQLcrSjlqWbSVfaS8S4kdSf4JKVmxj0tgemWEvBmhY3W
hWJrwv9XqU7ADN153b+QY76VAoymuhIRjfDnEMyiAwInEA/LYfqaNw7DGk0jmBTPMrgEukzKcnyb
g+sA9vHWQjYr31orNceZSJB09j2PR1/ruUFtbxXHsIU/Y9gpDMTSrNgbtxJNSbjd+cAuO0KDVqQB
zdhrezumplSYNucsFOvapS4OwRnQXnZBuakcwgGxpzT8eLmQwnlVI3B1UqTg+/MtHjnyZtudlnrE
BB193Q9qXBrP/12Zfaep39osvrSYKOfn6qZMbbnHnMhwy9VmqZ47OIDWgYmymRwT1qKrozEukEdI
MkT3uC/adIqmf06jsvitslZanwfB/yW/aWjBiqfAq42jXsnrkgvLr/U7U4CEeCZ2rYiABfXYMbJL
ABn9avzy8AQTCnNTwx4X5nRn1x/DJEMe7RtTVVa1fXAmoA23lLb6HRLZ4fojYBTTWoRJo57q752Y
efv0i1VxInc2tChAeMIzM/ywS9widNo6kwA5tvpXzHKoIOW7PCxVNilMoVlL5+AHsOuNyNBVykAe
gSYVYOCJyQgkjM9bceyPmBdIBZnGEpMhmjTwTWD43ApI/tf7GSrEUAHVpdfCIPXYWbm5oNGCHq2i
5ccBY/pZXkohLKwv+DgOetXm2JcPZDRfxBlLZeCg2HjnbONppG2OfQwNKj13PdF8Ek2nMxJ9ynVG
AbQEkhB7CkAz574mfGgtDMw+u9tBTJpAc+2OuhwtQ0Rn3z1ShpcbA7xvsAQ1G3E812DgUNuU7MNu
4uKmUGtaPWbG/KxgLdabgRwAULLa3W6udoKRfMibVYiw1mOuCNtYn0nHDKKk8GmrKhkciCN7eUkR
9IlQxeyZponpD67oWNwugnsdvfYfbRAwdW3bbt/0B/wqsZo2FXXl0GAqN0X7RcF5zXAA+FpcTq2X
QrCWji4RRzQ5ElwrPXdjb+WXugHszEF2zJPPSKp/WBUhjiBvrB4pWjjsIrgJ6zuBwhX52quUNVn3
D75z33U+QVFsBrt25IUH039oU49zeqRMJac0CLukpWkIqwrbkwzd6wdOQZFyEh04iyO1QNmwGiWA
8aEYbW4urKAiswr5XkHiOog7eM2OJNMVAqygxhGNl+ISt53aQhMqZECAYWDLF8KtbwxoVhF4pUPb
XXFWftggKOAD0VvFvxo0nozzjLQPD6BQivKJorGn87uJOfs3m6aFweUXU0tREBf8NVU34KlDN9TH
kgjaPpNgovZN3WpxsKFuOrjNqri2h0q7zxgvv1YYw/b+mT1njjY1toKXb5FcR8A4hsfveymC0E1+
M7cVSO5jOfLeSs/ej9GA7hqm19yHEenAxIb1AyG9fZl3z915M2cWKqZS1zpZHZO1N//dqXNAAkC2
JagrftL6xp+nqqmwjlP5gVEffXZr0CmnIFLb9R2X7fomXfV9xbLDRfDa26BYNK4BDxRVOSFlCUjT
hecSwZcUqF8kX9YpX3exU8KaTahBQT1lD0h26ce17Nihh+8ZWcoqBH25+8vDAoXj512KXnBwATcn
D4hlsA2SzYOPo6+5GJ8P1jAtxbPtTwja8CZArXVNFt7uaBWkX2C1V+ot21iVC6R4A6X42txcJeqW
yxW6Sl6V8pkNGhJiOAFSdFdWI/qHG5V/JrngrY9IfVRz9Vs5PNZbK800Tp9HIqvEcfaO327WL7sD
8QvJlPfDrJnY/6mu7aHWM7a5ybFujjgJv7e7d6kSbJ32QqXEEvrphf3Ovi5UeIvrFp7Mn0Hgoftb
kumFsPac2U+Is4JyK6zKJW61NT8hr5/Jdipo+e6KRp40s0CJIm+FgBqvWJgkVk/Ayd5mGknbtVF2
2bFnbNscp73Tefydp3FQOb8whdNzOU2xgELnTk+wFtQihwhCNSz9Hw+JenqrhaaWGD6rC7GMDhC7
djkR8F9dz1hEnlHG8ToE2kG7RqwvoSymrjPUETAES8fcuT7SFepnJgwE3/MaOQnTpWX6gmbMKwDU
wlJfotmusHBFI+xDBsC1RibqxOMwQfCnllwyYKXgewtjtO3u3BKtP0WKVHZq/tVOQDp3neQurkXN
6z/Y7hkQwZ4avBIhWklceMRq7WNy/Tl/YzgQ6bq337TEagRBcQwMDrMR1T1PdttbIfj6rfR6DKJ4
ejSP/NHX2piDLb5L290kbiXarwoGLsU3XeNUjjF3CSUloPFL/g0memCdOAMjgZQyuhX4dJcS09s3
ZnccCiUQjZ5nCsuUXFNP0JPD/L80Bbni0EDYlzA4hyyn9SsessXxTBsNRaA/YPGI8OzWoXMCK12i
rrr+8/tXFeepBV1mPuP+Vqp4Y1R4wF8TNmXUUJm/Xd67TcALh8yLGCUhP383TptcFwESpC2DmSxq
EIZ9Qyz2sVeTBV+vZxMVtzzbY6fOZkY2OISzDh1Of6PnaSHEnDT78pRfHVvkDY2QN3xDKxmaI/kt
1cSj7M2GAqxOnpB6yJlwhiJJ0gSZqF8Kx6P1+tj2uhOxNaD4NSKBw0el/BjBTeqLNa0h7e9CMDdx
GUTE44YDOset0+QnTtStgha9iNRXBHzutbK+iNyXNBGRN69kslV0o2gO6NDvTuxtyAqEZMVvohp3
nAqZWs4jEA91UC7JW6nfzS078L6SXMZ/Km6yRr1G7DwU7iFNUDL8KV7hqXsiE7GURpXclqsXdsDL
bV/hqDpAzHWkpGd4n7G10bsK3yrDmm6R+aGY6ZNy+aaERvvbGHCtEVHu0j29keiWJStt2WWpOs2U
k0QbpUWwIGcCebMSb+Yg7zAY6ODd6cACiTeN1ji/vidxIsuRIsZLbdpm1YoTsPLD7c2XLE5J1QVV
yUJfVncHcWws0gzegdbQsLHXQ7YApHQHPkG4na3o/Q+NhWmstUQbvDDW/YUBa4zbllmF/NzgkXNx
Y/c+hoWITSFhcwGnCq7aHwzN5TNjAG4yrfezd9d30IHVC0j3iDYr7HA7FJUq4rFIU0q248Q38m80
cYHxbmbA2tE9sA8J1gx6YISDxY06YnutLEYEa+1SwPAlrAO6Uf+CBymb4YT0YkoHdhkk3CBnVdwF
3H75WH/LNKmKkSWLb64nK+gTi2lojYqH7Ou7hj+p4Kpc1dZk5W0FxmRLOhxPMP+p6dhIKI8426xp
Fy3Qwur7EhVIxIezmnvHc8MQ8OtGn65QLF0iBE9GknCye1krDBiRd8nglQXBrq5YLQSwkpWCYGEd
7z91RbmLQld3MwngAMemepKa/R14kxLCrConeX1NAsIgu7ObEiigzsJMkFRsVgtH9VVlfZtFAvk6
UFhYZN2ILrNOC7QARYJx1MQqp0dKuibY0+3b1Zqv6kprRT9bBrf//BMUJ0sqfJzdRTnXJ9JLTj/L
anMAIdxQ5mRf+SXwG/Q4DeU+aPHFhSA6PzeBOCDR9dbTcSv5dF07baLXR+lALUaWqf0jKDaTmcwX
n/U0B7R/j0Qmto37due3hDJqWyg1EwKG6BDiqgds2KM48qjxC6Q5yCy/uBIGQez85CvHsXuRR7Fr
+kH8/NBBfviyevOwW+plQ+EgDZicRtxIggHliMBGvvaM4US8e37sMWpQZwD8jp2eezseuR6TC64S
qJ2EYY9QpLkW9a1/L3KCQuMgi16HOUGRgYMfHruFT7+B7GrofLNQS+G+PDnxqtoddl68jjS4b2XD
NjUC1UM91SD/zP1FxZjkMgdpsnGTJ3xaQPFzM6sXe8uB2OetGa+jHusxgZHmeartgNsTUCVs7UFW
1+oLm0zbOcQEdOdfNr1h5vVrTh4eDURsGTco6HRS9udqhBU0C+9elsfMWW2xxdWNWWERR7vkziXW
yiVjsMN7UB4LFpRCknWU/jfTz2p78wpcZthfA2LJvHCY2WTUVPtyKj+Pq9m1ebJSQ/RyvRWUANgP
EdGS+PGhzW3VDlSzovlQPZZn5KCgkybdvWy6gxRGBF5+QnH/LQPb7NdskQ0OLZNbJqs+Y+2yUQ5Z
/138UDVEOrWMSyWr95C7pd9doj49lGYyMC36GyYwaB60DtsI9o4IDmyMcYWPRKDcImkR/hoU7xAF
A72xbQCKXxlUPe7KB7/2AqL35H4Q8UScxBPUdQALg8iSSZ3SyYwoWGui/5eboyOpRSli182T2NKU
UcuoQcXaOFES8mNbNnrXi76NnWk8Fj7fkTquryljTeUEfTdMY7p/Kw6YUWpC+/DQMxZsXVZw3//K
a4IIec/6I1FjJAFuSHsfwGN5/ph7DnmyKJ2/nmaJQIV8SnihBiTHppMUWMhCbwD7t/7euLtBzQ37
D1fC7CyZHH1KKYKsXS+a3ab3WEIhb7Owc0hjGxKUTrpTKMTM4yc40dHPS3muQ1T0dctrK19Xcgii
aWpwDw9oXWM29VMHApnXGfqaM92i0dY2k7HUH65IN3XypLF+uWRSlodqVErDR/XIL+1lfUHJcWyC
1XDNdrGLZJL3UAXOVhrYaPbu7L9z/o/s7dv0o11kqBsAnI0XrX8L32IvfiqaXsSnZcKyHsShS3DZ
gct7rHIPgD/Hej+73/UkNgDFcEbuvbMeKQrvk9Qi4fivVHiTrNxXaZ/zcIJ5Y5COu23WXbU3GOd0
l1SHBHpfXhqmLsngc1+WapnxC87XCKAiQ3sIJia7nB39fldbtGb13SCYugrUG2cc8PSnBC05XGCo
Mo56qfI+NcpMLdZh7/MjuLYQUe4SdMV9uQj0301JW2aX+93pEcDpTCEg/vi084nAiCNn75ZkO38+
KV3KzuHiE3Fpi6+6RIWA9762wT8xsYgeGD6qsYjH0K2HxHAuhMaJ6IvIvnOlCVlQUsksaS151H8+
E8c+1Mw7+KJqkIzWB4escq+bDl7+RHlUGNTDxgKPhD9G2wO+9WTYg9hSeTqHIVQg4sTnJ9kx5md5
lp1e9aX5ik4dRlcwPfPXWyOtlyins7kP6btKgRM9fZuirXpRVWHQMvgUzV1zHrZfpZI1B4lya1FU
BPP4FT7Au9bG9DABmsz1qg9uO62Kbs372jR+lzUWU6/mrOy9mPETNs/J9D9Ypsno/LxycMJQ0+Cm
NdH6FJ8geCuneqJy8d3a9ELPmQu6he15goIN3VNU/qgk3maaW980ZBHwoky1R6tDRbc8/CtW2AG8
QCLhatn2FhW6A9oRds6iNThJWrO7D8tr6xsIdiGeD7NVuMC5s44Lt90sJZ4Mh+ky2cLjuAgatpyC
2opEekc+CY3FOt6lXW1b55xiyEXrP7CET1bXHnZxBeUajJ5o61C48PKQy5wjfwEsNtfc8ba7WI/P
PE1lCO/lMJqL3Z7oX/IWV28A4QfUID8rZ/sJOkkYLDsOgZX/yy8g7uKtrTS9sVMRLP2hy3ZrJQyD
KmNZCrg9+h5wlmsTfBsnvcvbGhjcKFZwGGZzlKwBM/amoUwnunOtzusjTBT1ViysSwOUuGeMJVhw
QflsQ/VfkpqSHPRqrZkMroA5HC+N+GbUpUX9b86QbA3qAmYRLRizyjfofDnPutG9TpJdB4TBh63n
lB+HPBb+cEqWVkY6VuvsOExL69HNRDS6Q1hfWLFHHGZDtEPfcVBHFg2AC10crNrQ8DN/aqB9claN
5PfVqnDaf7+5hIUjZD2gYM7iPKoYTfFf4osIVoQaWZPmyEWPLC6NQzD7HQuNMGkdtfioaCBdcjya
zGKVIqH2PH20gb3v8LRl5cHyJiQdbKlrJEsnorcVGJKXpu6MOzp6dyo+QFGXkElFEt1Ovzp2MYCB
reOoj4rEE70RlYT7xa4evNugqg6o3vkTzwH+lBTd/qwO5cMDy/d+XDgYk2sgjCn2hO8mQA4gsAn7
jNjlng8Vx4rYuP21FtNINIVYOd56yvGC+7av1eNpCk6NXFw0ylenswoP57YWGyuguGzgFO10+5km
9BKGQnYJF8BgkGYQbYgFZ2QUeOxcIm1CoMCF3CE11iiaE4Olvwb9HPoxOOsapdjzMF7CsmsirOmX
TLbLyEHzfXe6FZZmzqjQYmbFXP6OzC2uboPp/yGQe/OZAWUTUwLg/g04YPcqovghMtl3gAKrgjCU
/EkaMxG6TcIHA/XiCpXkl9mWdvA64ml1o9UXlbsmeSyWqfEVUVjWKnx/27BjZhuzL7sFVq58XPGZ
UmxzoF+lfz+g6BDwABdI8Rol6qao21rRQZWNCUjhxrQDMDELFKrvVxcQyMGQorJ+0V6lZfYa5YM/
Elkj4b0h2uWiwyn/6DLdxiLEN7NUdelh+fGQ5k8nCET4C3c/qwzJLXds0l9e7HwiqHB8YOO5GLEO
N4daBDUj5eSX3IB+iv0Vi+LZ4IrwigGmW8SZyeeQsKBOdsYGn9Jcb7Efde0HlFfmbID03bAE3QPs
hOh7SOUiwj56+ekRFTXS7rKzP1rLLEpMVrNPcj4qgUe4Sg5SYh+etjzXFBg8yc6TN653AWeZgiW8
Y1bFWDErnoZuUlZ4K2IzDLaUy8/QHoH8rk2q1jC5znnR47pa4xAXmK3sSyoqhiYiJN0uKTyvziIy
idy0BYcJQWYsWyAHhsynCQyxThjsDWUEejs/GXFbHV3A/8eB2EJVFJCgtEPSa8dF0lPN1SgJVjR2
leXlq1nb8LXkYvzxOtWnbOKvGvuVuHinfx0i/lVoFvOAS9jOO2BXPo6W/kJH/GE0rp9XgWJO5kmv
fo6/ns3/22ZnV4ddNbZl/MuUPrb0AYVXgRAIUDkhxsXzjZC14Ia0qRWqj6EwCbEL7+Nh2LIdgQCR
ySEjesSh+Kqg3OCZeh/+0vDhA4RSquqvR0BYzr75IJqlMzKEMhXmlOkmo94wgR+Os/z2FM/sZ1zC
8O3hhGmn0JhLEadkVahZYxenjILGVng3tzNUlKCclpIKwtU64wbFq+NCkjRZgsY8YwuSc1avvV7u
lnFblzB7aGFHNoKX0mGEtF8a+EYuZpiZ/GurZCvwgMo9XWtvykKay8Hqzhy28NBWb1n7Ud7wHoMz
z56h9xcG4dNKDViFjj4wt28TLmMt6msV0Bj7WCDBSoqDEe77CUNYBq6bmr20kREOghXEjimlYgGa
sZ9+MaVFfBNVlwuywJyuDV84Xsez63Db6eDrc/s+vd9RcrG+DboKTWY2CZB9IoEwP4sXEMuFFI2W
PS9PqP/vKRTQRk3xRAAZDhH0QxbbvD7om4fMllzfeX9dGtVlt9xrziS4G9sbGeIvSxanFDRq91hQ
QxE8kVZJTenfK2cYk6bamN/ulTZKJ9rSCR9DXrywq553TMwYvACDfsWhCGALiGXQFR2/uxC43wS0
c5FGqrSgD0GmheAT5rvyfpqOik7N9yfAPb5sWdncDhd+MVD5ggkt9Lk5gPFM17+laUUKTr+buwUI
J89QgQnqGb1U5iubArgu9fMiC8tdkiO2IlCGy5wEZj5voE/FOvYYY5xHpouBgHEx6Hcf9YKRgwfC
CqxYJAIYGejxMzrOM/RnOxcLNxptrgVpm4R7aclcayQnKPPT3SdxY43Z+PV7jBugcd7U754KmqeC
YmaT5XehS4pkxiTwKpJdOY36NRVOQxc/fkINDpv+JmpwTUMApnHi3y3V09UZjasEmhBjIT8GdsWA
fvWqyCcQADfx1XXCEeJnaegIQwb6RrwhWJpKNHxZVCl+uW7HtHAO3XKk/6kaqBSo8uVHEhoTd9Ez
SJZCan7XVV2zzLtJ/4W62IWM+67GQzWVYVzFDtrEq2Gq9AVglPihhbk5FS5kxhJ0M4rEbRhCepvq
QQTQyWkSxG05kUP++supkDJidzyZsfL9rJSP6kLgiyPt81CfWjy8OSdA5MEdAkMYXx1Q/yoJykY5
7UrKz0MbYUsffJqQk5+FfLit86FAQCu9PA2Yye1vyKTE1IT8M7F1H+RVRgzKgbaYH8xIYsTdtU4F
5QyRcmdNlmND4o20WyhCj/0pCYQ3JekByjx9CS2u7BINu3kBcA0KjS5v4YXJosOiooRmPxJc3KpL
fYHqAHlOL9xR3EUga5YuNSZ++YUnO1X5SJIMMyYl9bDOU/fsXel/owvt3sRiGCmHj6BCX00ZsJdb
1pfinGRoIJs8gnNBsP00xS3VwPbPhGc3vl3Wb1D5vRRNr5H+jp4EGDHZ0nVjoUEeV3+h6DRMyLNG
yEpFJFD055vXcpRYvOXrhvcTr8uQFtsk00Lsd7SB8gy8tfh1QZVNK+1N4ILzLcX0bXVS1zMaCE2k
2mLo66t1kn1ONmkJ/p4cmm1ddt2hB01vqGERQRZDDIGp8QHg/cg7ZnyIVQwdwT/CHmR7G1ENbohZ
sQc2lcPeTq3uRjGhdBUe/hwewR+LMGIT4Or6NrSN74LVjlPEYg/9gw7+agVlXaTmArSuuagLFlX+
/6fxxP3QTk97QG+IBMqr+giztwD8TIkJbrPUMK6sOYNB7vp4kVFR5Wjxj6S14msJeo00GEsZa3dQ
q8g8xtGgnlNaalBNVX63/hp5DQqlq4+sytypXotnyGxCoG2eAi9+hc3tsXF04lm+seAvfaA0U3xH
2AVSxtq02h6MXVforFZhshWsSMwlP3z/wJLM2AJ+fyIOt+fz0tnECgXhJxmyyzM5Hs1YmezmOpY2
mKOnTs1FcMsCN84LFsBngS26FTRN1l1O9DG7ppy/gzYGAhqlt+aDWtPliGmKrek3XWUJn+to3bAm
tHSLZcvfTD7C7DeEDD/6VnKDtJRlOYh0HB4b8BTDTCJLdWFNNuwrJhnloPH6JghLIhprrj1eCM/L
XesQpuoWRzYAyQoRh3GzPJHTVydmutGhMtxodXQ6xZw9eeNsCp5teJ1JcmigFtH3ZEVD+/lKYJiX
sxF66kL0DJXVwz7afm7yPqxl30YyVO9xOgcBpWsOG0U8M8/A0R1pkYj0YUAOkFfxjQ2QrZI3fbbD
VeTuFfS3zhHmFV5D9oPkDn326zmwWMfeYWFYec4emQUk+VMveGEiwO2udXBCNi831KVXff7nJXHI
1S7kNZNmU2z74xK3yCALGcr+j2U2cxmC4QnCapK/N4JTFKTQWXFxessc5RzI1tSUg0Yv5QmOo7En
OZDdRiY8UI2BOkJR8PvouCxX5hGt4SVwDWyquM8THo9eCw+Ci3zxhpTaO3ahKHmZUm9zsbfBQAjn
pF9PGG80IHaHeS0+YD3m0OriBrgRZepVQdjsZq5aJs1kYwUM1K2RW2S4LNIZg+q2LXAK+38anl7F
THD4zlLqmgiXoBtpsH/5kuA+QFoL3dJQJNJoHjt9SahDwOhplLFYVUwcSP4MK0B09mwQH9QDz8XC
7VNVD6d2qOjkjpEnOosPPZdxJmrjs3GkupEzPJu2EpU+svI9hPwXik00+iqkWYjw1fPMDFZu8l7a
TNzIRhCnAJ0bCdEsCQQfx5YXI7ohsDSvm7FpWpI4zJHDdbxN1EKNtq7k2/tpWrwx/Q4nxE9N8+Ci
uiWHDukHwMRWa70Y5KFQhJRWo9ccuVPHkaH8TSY6KIjHqjE5CydARoOWlCI5EiXZP5CH6dVBru5o
SxP0JrMc9b61NxSeBJJxgBgGsuL3ZR+pL631yIXoR3iCnq44obcI1AkfC0fKPSr6WggeOzrDK80d
eOB3z6LNKTUtDF8WTzcOcVvAiQAD+BlBNyf3XvtT05ZnNF4RN9zIR5IYjUnN2vSiCFdNkmFs5uMq
LmBIDlL2ZzKwNEu0POdx0CSC+AcgwLN9Zg3jc93R432F60EGyLCTMyN8F5zCYjlvjALtHLxQ/K+F
CNjoH/s5W12BndUWlF4Q+3OvEOr5/MJ1TnS0ar29ruiKIxmKoh2zPVE2UryHe3IAMJEI85zaZvWU
HfMjjuSSAhT7GAaKhMKGbSdSv5gWOGpSzSnAwBskEoWwWxG7Ou9qLRE2XsxDaul3mHhvfj6yb4DV
MumaNZfgN8DteooTHeWM59AAJ4mZZKeARge74vAlS170mFML1IiwhUScuL9lwxgdbOTcxd4doz/J
6SeU/+QlKgeJ8IObjmFQWjLG951Y8j+eii5PC0GMrjmRQ9vDZO4COvBZ6Shm2+HH6uD5hfh7brxA
1suMAaRO+XdPzFTQbdW1gbsQATutUZsFOsRdxnDohMea8PCLEZuIdEtt7OBCRjlweTdnD85bDm39
/QUIRr9XyrWTu1pQZNc4RdsY+n2JryKGTguHx7HoEkmcoJRp3TefZi7YpmVq4BWxrXqG9gFtPo/K
6yG2fsVpejteEexjaSqZFy4rKK/f+Rs+wihsJIZYtRJXeE1JR7ILa5Of1HSTPdSj3tNMGtQ9u6kt
f23F254o/MRshzYKZpixNe5ExStRyeGF0yLlteRJT1lO0XRNe3sQ5UU5q/NsX8KXXAdvwrYpxiri
bSCP39qXOLFZnXR2c3F1l7SbQkJODq8DDjHW9nHXG3v1fdVI+C5pgsFxmA+Y6JgdKV6cFkL9/5aH
KnRPIDyHPKtJ+xf/JoTtD0CEkxcr26NQ1LGgYAGAB/bw4t1zFOquKNePuKafGodQXeBikaHghrMh
mvD0hJJI9oCJycvdBthEEjng+4f9P+MxeyKdQGi9lm81AKRgBTNIaqQmqy4a6P+/eXnqPHV5t7Ja
wVIRmjF1n05Q5Vl0o4zXic18RAQe72kHUQhqCdFnRF/ZK6kVltnABPTKS75QIt6c1Iruh+oW4IAm
EvM6TiDkQDER6E/amllPIPAacU74InD062KRdcrGGfX4mWMrkHRb1DewNgRyA7B5O6rMifH+fMPy
4HmSVoaqpspoFlwZe00rwsrkY8xud4c7I7YpaqnVL+dhj1PBxJnkWYdGR847q/Ti/anq5z/JnYRw
uVtij4zJGhwkMPyOLzYAOQW/46yEC7kcw/PvHD46vQwTyglfDy5T0wKGiUtM0a98QCfnBceX0U5B
79/OoIkMv69nBw5jXnutNZ/G8SeDABdYdDvK0qVO8erJmExUcznN1/8uuwxCQvmBxDszf7svSNXI
monY0c/UujLb1gA2rVSsqsbnAwagFv7fmHF4XlD4O4pU1nQT1dLrLUK/8Jin70HZrmgURhUnbMQY
j19OSsq1tGRm3+3BEoDbWDbAyy4YANtjoRXGEXMx6lD5HCP6d4FMlXRFdwVOG6Cn5FL73ah+jZyu
81yHu3v5h1O9XHXWgMMkCD8pPqjHDcta0ZCngfK4ErF2Tn+dtRlhwuAvlSODlzAGvP2rU5P86Z1k
wWE5cCEKe85r90+MxVS4Z47dz1w8/Jnw5E7tgsPj7o9YKNj1JJlOR7s6GozslkCIw0bJ1L/6r7IF
4h5X96F0ERGkxHLh53ModttILxnmUytrWuRY3y2/8j2TvSonFsIN9gDz/ncoz3/D24ZU6jeAGupG
TxC7rAPaesaRplR7mALYJrsubcHqedAYXcHOLZ6xZ8Xr/q7NMR1L8V4kW6hnFeyBJRKQGevQQRCB
EsYDxPcU776Qewfqh8JE10AtZjqzKEYkfl5CjRMMkD5RS4C3CZhT6zBLh/vHYnPDCLqTcoXF09ae
KbXGt/wmFMi4GKmRdOtXyh6Un/kn4UyVvrbmQCMLyGV+o0nDicIofcHxYCDjZnt2YEDLRdtlsqR3
IFZpome5OTLJ26ekw+gGITpZzMeClTuEmE2eCPUenME2djVIQUCuskUBSnDlo9O9fB90RPEU5qLU
XX3khMCy8WIJDn3ZUyAdO3b9EsS89B6do/VPgtzG+8Bco6cGv6eWTy6nynU1CSpirxlI+itI8PsW
R8v0tvRPYIT5WqqW6S/HT5/6QHdIhvCYGV1tQpfKGHk697Ih5CvBTZW/3td0gNCbcG6iihDg3eIU
28TfklwgTXd7rkomx//CWx4+uoR0+N0S/YYSIbvUj4pfynKB9iRoUTGb5OYOeG82g5bP+TWD/lYE
flBhV6QqYCmlBxYrItgq7AsN0FdWg5Ple0ZgxC9jSF9/RWWofowf8xFr9ejcnFd8dDeKI44zpVti
zYyR4+Yugl1HSPy7gGOkENlxsc9sR580EcLut/uvW3lJj9D3L295a6P9CCUGuAzsJinDd4ff0pYZ
Nqrw05ilvmCFy15D7ulG/o8+X2BfFTaE2zZH/0fPl/tc0JR6vXDbsxtCQVfRZ/RYZzD9lf8Jp4Ew
yAIH5lLl1sa8W9BYBx2k6rijllIdXZQM4VibKhPo5Xtyi2nltWrFOp+V0cxK4dKlvA/IBa/xplNR
XRgHxxOM1VuaxNvESTca8vh/zJynod8JjxPyveorUxZ0QIdf3XyishrUui+4R1TSkoSBJgVY2tz4
xVsezD5Y6CK6dFSyR+aGdLU35c7f5L2MdQOeFbMNJIftxsWgcma1BoWV1wplRIE343L/HoBnIbFs
Dn71Sj1jmjumAwexzfQ8UYLDM/pr6Jip8jmcMUnAuk8gFNdesw7YXazfZCiNjCMqDQaReCG6Hi53
g5ckgbALC5XdZNnX48OwkCM4WvlsYjf0YrqmzNoxIY6IGJJMit/24NPzDzwcdGGdUKrmeSde4L11
/pF8aP8nuw0rPMc01HO0pq4MRbtPMY2NLrekAAuMa2kkAPNiQS1BUHxAS+Dsm31MKiMOxJQSLggJ
6jghzkWQQ48cZ3AZIA0g9ZHoElrKZwpf60/arp/xemfLtjCu7aa2szzIhXxUNGH0I2uzLL6kwMf1
UiOQ/veh8zB/9qkoKqUxUlAlvZmFuPsAaL7ntD4kzffVNmwtj1i07Hkmx4i0iLnLRUo/teMCakbr
tg2JE/aQxFJoOrrkxZpKCsZTlgyxjFYshbCUPJJJo4F0Y2WWu5ShTsI0Eqswxl/xgWhr/ZxHmG+3
gHtfb6dOqT82XvyOad3GYHCElCnM4xzOv4wrlaaBYwY0oMy1NtrfBygoIXCHDgjBEEgrVZxdKsm/
0LPzo8ukQaMjJGhmjDDkNCVCHA10PWNe7aOIDMKFS2Db83KFWTIjs+ueWmUpJxlJrK2l2WZxtItJ
I7soy9zEQwnbqNkxbqw262Yj6FJO7FrKGGinFjn/htV3ECB/jTyzgPHQ8kyF4kKxA37UB5dywfOT
vB/2YudykwD9x2T1087Ee+cXbh4o37/h4W1AWVMHLKKgQI837Cwl6Hi/8lPqbFQhuztDYa9dqwOt
D5vZtP30WnznSWN7LFwLjoVlYQ4BHivbFbm8V/Mzek9QwxSVmRPGMTRMtmdzLdcT7cRkVFa6a1dj
sy5wieUSXDnexee7xNH4rG1kZF4M/GZnCfijSp1CQ/sHQe9todXOFOa8RkfdF1Jpzt6tY+owmxma
k0FVC8vMCY4uUNQcTlz8Ua9PuZuy9Jy1sKVl5vm1UCzYcG9Lm405NcteD75k7BneiBqoV2VFX79V
vF3R6DY+2rpmuRrVZmKXqBcO7Ee3pConiKfmAW6vfleJvuMEO0iNOAA6V+y46Xwb+oPdys6fNa6x
BAcnnfdVq/hVdzlL/Ertl3tkUaBmy9F7nmdMQDsjNaE2VmxJlhi82XD0EgIaGm7oswD3OqU5hEik
C3z06T5ZnACIIK/qsX523qKpIL69GTH1PbToZ/uJ+mxmAzk8Uylw3iVi21GWLwAQrTl1tapWHX4E
8A57jhr9U4cWYGJiTPBBSunXhlDVHKrFxn0WgH6kiyXtPAibIBpLslUzAg7V+eIznAc2OOav0DQh
9GEVV9gVHYjnEBJUTDbsBgtInCxVQkBfylddn49Gw9EcegJoo/Q06MFkIYHXERj81PSUa2rGO21j
XPVPOB6omMIbBn05hVxviCmOztLPW5kO1mfOQvE2lxs/ugGJVJcn9XDTgcADQ1ljNC2/SC26rr7P
8dx9xAaDXole01+7XziZn8nQts48G0hiF7BbnnehRw20I3o4IFaxNyolowfT0DlQ7bPNIRTJpG/a
pn4HeGy6Cx5Q+Bzjh2Ona1xIWShsT5s40oxv1Y8tKzxdG0h1rIahxLqpsdQuHG2TepM4N+vLX3jn
kawnTazvpe0MWNCTUOwtNXVOYngrj7Wb7F/uVjJKBB8fy7xAPFvXi+OsMFLmetzBtYXXjDRYRgPc
qzMBRUPDMoiCBJ/jh45nd031UW///LMS8IW7Ym60VL+NwKrOyqQJ775a6c5oRtDGJ6DrX/Sc4f1w
C7il7XaGjnCCItopjs5sWianpS5LKVB3FKnhKxR1Kw41vBJ5HPQWB6681ouWFpnNQLfujg0hPXqe
l5mVZEREyejJzC/a3lnhlMuPvXdLnQ/QIiW1DFhKDdtdMM051qlv2V9rQJM63qMjhFeZByNxk92a
j6AtgM+U8Vxkwa3HoHLZv1bOnQngBzLLodHZWeA+OSC5l0uEQYVnxfxx7UDMNI/A3Unpc6mySpFs
NBQ1WCgiA9xTVSYXatbaTw8ZwAZP2dIqyJtiLvAvqQoQ3Yqz6I14n+feowkO8CUtlvhQQhU6Wcvw
We6CtmtJuN/a5GPrbojzKrrXMBTKoiVVAao5uNGhEzhb8DwYguuTnrpI/6b1vwRXnpI6vlxHzLJp
1lafsuz0bsEJZ1wjc+I2rHg4fkzkq3RLdBCELBrA63PYVSnb/qFE3VAQMJj5ps6kArCGpvgekOa+
QZwtBU11B8Pnn7iq89gAi6Y2vq15dD2UsCyit+6YbYdGthhzyH53n4Q/8H/xzdZhyd2FK7FYDZye
RGp2hgRox4r4741gGBY3rAf1ArYpX5eg4pr7PgZ/Ve9Rb/6EUTsz3GiTYewwBGB2ploVqdqBWZx+
EUhxuA90ud0ENbW0FwJXkdDQr3znDGoVAZvliXFrB4eOZTMoAcsrWh5AgoEeU6bV8ruLSJzp8za5
bl4Wt2Wa4Mzx2TH3WFT1y2sxRDkeEBBpq54Ae9osby3hBshkmMtXajM4LnVI63AQxKJU4w90hC9P
h9mL9qWdv3V+L6sTpadWkEH8/uJR7n6WWKjDzjZ0+zLsDvUymyoQyshtmA60U1FRme3QUAEhprYj
+XL0C5cDkRsoWKDEhsdeSbvXfAVxb3vco6h7e4wU1PikAi/TZdb6LOQGkI0XCEuHZhHEazAlPSzx
amhcxX1Y+CKGZ8tb1UPR34DlvWHiF97pefppD/fdeHvY6SGftz8lrV2Ba3T3mQ15QLQ+d+4rT63U
VEM3GA9l58Yvqcm2x2z2NJhO9e5RSAFECwZ4mIQ4elZF218V1UNJJ9ckALJnqRbo+2FTDggyyyEq
a3Ka9pO0fG50DYu/rkXdX4BlfY030dExcEvjwOgSGfMN5qv4WpZLmCwlG0hRgK8IOlyczOAJxkWb
Vf+upZH0P0vXVlU7809egan4QDMhq3875BUU39KoeBA7FU+eGk+DI2GjdDEpMkcsXDktUvzJrQdo
lMgypa8wq3/JpSwhrgzKHPKWKlOZcYLR1JQ+4B/huUv4NLXYqKMOqAVSb2I9TQJBtkZr/LPTs1xA
64VGg2+HIxAHbE6cuc+KGOvcKBCOql4FSfBYnttdo0EXg6YNvlXFAKSZSK+MWV2eU2WJnGox7hjo
bgYXnJWCmLS2h8IwGURrLm02Cwew/dAPIkmS+An4jyNot4DTHn25Xt18FwsfxlfbhUJJWVdMHpkr
kHyngaTtJPb0XEJQeM2+ii5uJxTJYJ+OU52/9CsXwUHqywwpdv34mHvCl46V4Cf9Llx/q9v6+NsT
YcOwmWqibAc59N0Ixn97xEmy/+l/CcBE041zTOsv3ArE5c9+SG6Pk9ToFRWBVaRkOBWGIKEYLefp
aMXN4MGqN5AoGQifCt0YvPwJ+iqzChq8U0tn8ElcgO+s2zV/hGf0YfgGSFL6S4F0gw5gUqZxvFdG
7KxkeQvMLmRX1+DxI2/64K/jsdm2E4higaHWTPBITmzPWiYY+gj2nF3gP2w8cO/w2wJllf8M434k
F3kYCMWl25KqPSLccv5r1cWmsqgDpL/2fM6Zgi+45Chn6jaP2EHoUUC9RIq67XpONsFGBSmaY4id
QHyMjOz5/6NkuryD1D+/+WPoHryR/cJzi/mCkY7mMgjGJfpSWex03muC7GjbN5VGkY70n3IlrE4j
0WdT0/TYLgORItNHiLriV8K/Npbbandg8hvMTYYVN8YY9c4oSMqkrfPAJIwgiJor82zP8DnIu5Hc
tjp5x11woU3snp8nbfd1OGWHIJ9IBl8qBTHTc1PPgZHPd+R8N8ndEvyRs6SeLfK3GQYpNTEm4Ka3
aLG/TPjOfaGwHAR/3cy8/HZyKzrjGtBZQdgeRMyCxYQhWNFgvwqxw0TpI5ioHACaWollYAr+jztq
w4qF8AxZ9e/ftQlvdl6rpZDHMOb5+eqUL3oUctvx60hgzd1OGu8DBjWqRcSN0M/YyOIzNanmzwlR
26fWfMLB6jgAkFDcO7b0A54bj3x5ceeO+O23jsdhhfGqa0pfBE27vmjHbupwOvm36Ipp6phFHtKG
7BpDpeJ9a/E4H4KmIak0/1XEgG0lh87W7VLWAw7rQk9GPJPXOkPBB+vFUfD25RMiLWYrxNl5Z0Ay
exa+4zIJ9LrKu/5XxYb91UKVJVrJ0VdaLcigQPn33ovLzHy4FKutNhwwRBLqsOhf9d/klDx5HlbB
M1V99fRCp2XN/lVKTrVfgVuYLFufmZU7bhBfvPTQkkBEV1NYgHRk71D6ugiYlAND0UpzCeS+uzdq
khY6xZqTz7fVNFnUO0eF5Ax5pYvO80aMxjbGpYkYx82yJaKLJDLhcI+ihvOGNcnEHB3caLAjccZm
utJgItQlSltGw0lCrEW/X0ERDO8W0N5OwMvfM87+tmt7adJyw00QEvm0sG6+2zHD43eConQfN3aN
r4tE/MjF6ZI/uYutBn9IiR8ELvlmASqu9/hdG/myNjGHWa2EyfkSGupddmetDcsRZjckKqhEiLCW
cezPFvj+ubWCut8kCxYePUqSM6Yg46lS12c2tUcR2Quytp6bS1CRwMEb3AUSoyDzMkHDgTJ5U9DD
xjcYBoqptHZac3KEiB+bfFwQ0N8fl3L2IieFHyvj7IiiWuAMdOCYsiTu91QskzHBIBKiMMh1Nlxi
a63GuQuU9WyX8seLavuha63zjsazpKUXSD9vWb9nsSUZ2xCi/Y54TOSCQaVMRNf99u/V1cd5mmZH
U092kOkpph+ayRVX7/wEz1cZcSQTTjNBUagVMbu9OviyFS/9K4S9V6Gss8EFd5qglLG5sXdU3EWZ
s6OMCoyxTjb5WH2sXcNr88ButE25DLY302Gbk85COUDnbd23jwwO+3Byl9qb0HrQqKGdzmfVas5p
aY8tXpw43/ucnetKKbKHjZtZsQApUuXSTLJ070zBd6CRe1U13HAcgjEXR3Db7UqFkS4M0/W7PdBy
lkSkLDkYLrHYtWoen/6VnbtTUli+3yJtsdRyYUCfrsbfLv+6/x+J4Z3HLBW2uS6hHLpczJUZrYJt
iuCVpBMCpL5OE0KaJIZEVZto49TT0WRBPXHjtxYXtnpmSwcpHXkC8LEqgCU8yBkVV9+NzX2EgwS8
6byHMYvRzViCK/oAflya3UeZ7xTk1tMSMuu1XZ5LKEgCVRIF0TUg2c5/I8LNBsduc2RPWxGrbBWM
WLy4G9u6Y2IG0TdWmhLV2LBouXADxmXiI5yHmeC3Q3ZlIrnb/27xA3NRVdrND5g85uiWnQ1oldRC
8xYCMVr7AZ1etRVMH8rtjD9JVhDxSOU10Z79PnenE9FTredg8mkcaYSLeHHESYJ85uFv6HVAFrY2
+NkNB7p+lpx+BvHlpLWjr+eI/Ieu9Sfpl/DVACzhx/u7SGzvIW8pW2necv5KPIwKmxotg0Sp1w+h
i2F8BbEe/c20TnK9gwqGb1h07YPZZrpABlczIAZ5dyWpZa8KZOv/KP/bGA3Tjvq07RkXzr2hYsTn
fM1sUGDdWk43xVx8eqBkTIPXs/WHaZDXwkO/Bw3n79AZXyzF/VpYka6blli000y5iLQdYN2Aq4KS
HjhzG79VGoZfmOWis0dEaC/DM5rM519cdkyz6IKbpee3L3uy/Jk0rVz21q9A6B1i2DwPx4yytuTi
9pG5XGzM+yMimU+2T7B1zFqBbPoWTw6VG2VFgITHLA8ytc1+rBiNy+WwKDN55IJOY5jfK4aa4ftE
jSUcNuIaD6PBjW7ZtmYcY0K1Tg/Oc9/e80SP1HVj4b6+Xa6q6k7/1tDKcM0nitMBHYhFJk466dAY
OphyGqAQZZB9ddiW2LazF0tFz99v/F8rV7g8MVw8FknjTDK7ppgXZDmYhHLxUC/lHSyghr3wiidN
jCzQOE7H0dFYxVvB+oXIgheWfx3Ar5W7Qfej7hN/X3k+ZQFU7gGAUKtAj2LPRKL6non0nereJpww
cgaDGSdVYblBSGLLoB1lIRDfF2VZFoL7nT4WB5mXXNy4qILNQ9l6MsPinJtOc+eAa/zjWMLdfJ99
QP0B+HcdRU/lPcAGjEXT7vBnXTaJJr0P63XCQkJf3brIzbV/j/bcLCa/qQqaNAT5YhFP9aa4Zozd
zqJMmWo/yktcA0t1qVagCI9MsuXGWOnKbqiUuyq2lv2KU3BS3bwLUMsEJ9p7YGRiERoXm/8WANvc
Grmr2Zzrhlwljhg6+toQBBQxNdKhhIugfObE+T5cgHfPI/VqCOMZI30GVTUEWuSbQZJTsroPH++M
3ge0P0KMxlAlvnWekbMqHbTKL8NXKwgA5Az0jLLlktvl+gFIkyFB6yy33LnUv3+Uc3E/6NNHmb99
JSUFSQG+fqLsL+cvEi/4mGbd4h0CD1RsKsd2MLev9vRdxGoKaKOUOQyJxF526hH3Nz1wo7A2K4tc
GhOgebD3XLafVD5la6hcBWCz3miQ8BpeT6vKMoM8CF5ROn8Gqz4WZXlc7VE70auF3tyXiIGok8Az
ioPMeLYa+pBNRBUqX6WEdvxGKrGr4Oz7cSCqRFA0NNERXNmUoiZsZ5FpD5MKXg4fAmAN86FOzdie
1PTd2h9xurGLZALvCk6WkXQT7nstSNa+JZyaFPRxb524DWNyHS4AAQVjCxTN/2t/S6uDq1IKZfVN
/aeyBZZvlUvnog/rWiFzd5EkKRnsFy/dEjAOZB5FDq48YGdl1UJTbEp6cTJnJ1/NiVylC19WQBRF
TZQ8TBOrtULmxz7cfw/lR4q9hVqISkbjD2g+mhK6Y+BkksenBw8mVB3Bb8dbktGgKNKxvlJtqUgY
gI1n8BbSgPjw1MSAJG3wHUMdwJLuVvdNyaIPOYzKtMH+Lrpi7ZATge3Fie2EQDmA2MrfknGeQBA6
IRN7EfHmG8WvzbWKQnGL8etX5buvh6ItVObS1EsAuOztF4LG03Z5YdV5UHA8FI6DmYItUowclIko
6hDr0pvAD8UgBdShC3XqOYjjRV/q4QqKbPAR3xrUqRKXGdniuSovVabjt6j9pnJ/+/4LXIWqXFIn
tEaIq6UJpBt6gTy/kQF8enxf8/Za6FedFm1S0HzWcFEanmMtWLMfCkWKsBt1B+8OQnZLNELy1F7F
MxHSgzdvkju5ivolNrJ6ogBKcUhMFmMHoF5tJ3jo1KN0zzo74wknqITd6nAqvuuvXBZSQADLtIDw
J8WLM5NlEbnx+jNSvrFwcl4reMEnuqjZP/vqPWSuNvllmI9U75RX1epuvBqd9x9+f1okDXLxXMMq
YQmDQHZSmFIvbawX/VkwVqAOcuK0D7JEUNrDexczivl7rDyJ/ZXTwpjCyiH/orJw0X8NpV39TlSF
izi4AxnoVTNaI/Jyy7S+V8tV3H6i8Uo4GGfdlgZkl2dM5ioL5RPdOFn2cDHXsworAFNNGVlULsqm
Wb2AwtC9J3w86GFW/i3OnpEuB1WMB02Y9SORx1IuKOxAaK5JOouJlIxyUdQBe3Urtf5UZwzX01kW
PC6Q8y5r7psBJcQ/gyot7q7teu+XCmRN72Z4XbeD2H+aHjPOMfw4/mMv1DYa943l6LAsNvxbN8HL
errOEfnsaXo1BKNw7tkmCLANSHwHSfTzcxqjsZXo8FMbRmXbGxwLf+tOyr+ps2GZWCJW+4N+cCCq
IA+Bp43xhzWAY7WAPipp1i9dz6guCBhleTwFeD7cf440h9ypKTDP9zFUcfbYkcQHgpaSS4a45wlx
izetuSuHPR/vyhdffVIc67o8TWjzqhGL/Aq+CC1d8qPEYzyr87hh6LEye8QSM3K/Gz/xMtCm9AdC
PkJJCmJouPDNbiMYVHrpuMA/TlD7Juao0+N1NXhr912CCCm2ORRJLb71IDFmOgfncMrx6uoN/CPb
w7y57XT0HlxGgQRapWDGVSimMqzcsv9BmI29TphsmIVStf3V5eo2Z//mEFy0gJx4BwfNoq/W21tr
AVpFDArTSzL8s+rDaIqu6hPPy4f/P8NS/7QeCAq6QRE+Qel80UNB/4+hQdhVBhuWyeBU7KFb0fwb
dZAqgO8+1ZvlvTvF63LVLzo7hHk6qqxUO9SAjNEEf4XhuSzWk6FWU7ymO9QSYYwjdln6ui9X3kkB
Pnfgn7Q6WH7V8tOpUdl42MZTJyxFshTp0WgFVHO8LR+YVEBopnT5sArdlV8IXr+Z/sezxWaSU8tz
ZXQ7olvdt2/lxScfj0AXjb3OVVqeh86IvEoDN6IPNh/NfcJdSxJYDBml4fvKShc5GLZqy7tcPtgY
RXBPh1ix6Ln4f8vbBnQ2RP7sOEysu2OcR/QloZjwmAxTap4AZaUtVOseyxvSBHpWTzPaKXt1sUex
hiHoaH62hNcmPERzfaHJzMUU/VaprURU0hnjW7Y1jDAN24SQmzhcAVuqRvqyRLwKCHwY8pm5S/eU
7DpaWu3sfUZK9M2ZwKSNKlqWp+awEFlf+20CQHmp61V+q6JCBfpEf9VyrSl9QTO/R2ZWXChLZkh2
ZjyZ/e3JLQXQFdS3w1Ueu4eotDosMq9G1Wo+XSnBlcV/Rg9z3JZDWp/O57Fz6ORzSmc11f1vvCjr
QJ89MXbKWcXJBSXROOeBqn5ebsXJsotrVsZw8UNNaxawVHnw3JRFiMMOBnsz6D4FFJPdufpqWr7u
jGcPJ8Xc9HkW92cOI0ssWkDhuvM2xnK0oKS5ZkwRGbF1Rkkh/oFc2qRxplStPrkSugwKd/M/IdNi
nlQY4Ew8LqP2P9MYNJjW1RczgWAc6a6NosHvR8v+659YMlUpa7Uk5kq1wALd+sXiv8574DVCksY6
vwQ9GT79tP/D6MLDAN6J98kGA0zqv+vmdo7o6kMinB+FnOZBzs1b92LJ35wCTaTWbKQznz9xNhpN
F6jvtFWz2S6W171Fth46WNebFQyl2l3IezpcEku//SEIKin5jnLIUsyW+T9wpE0NBywqOvx9xMlc
TFxNjNDQWpjyuspvoOCtKCzjHENsR6vIS9TgCSH5wIRnCNlyhUVue5KsopVdEJp5qfrFri0uvf30
Usplv2vxQiJ78TACmLflGDuut83HaRaD5kskCz3vxqqKmSUUbzEhWr/vtXVkxtkkPG0Z1kWznPOR
zi+kJpsSryMEsxf8mBdHI5qjpkXzniUQcGR2O9rFIK4YCrJilofCF7eI1uRH8sVgWgjWcCt2vAUx
lNFAaJAkyoSys6GjuteY+zwE4kUR5X2H7YawQBwQN1QlMZbR3SRihDujbdEGP2CpyLFifdneE01I
TDpTUrkKcOwhJPtTSPXxeAgXJItPA1hWkBUg34QX2FSGGDC1v0kvl7bkCyj6HP+hy9zIarhTezpE
tz3jrQO4bGgEHZrVWYYRwf6CQYB0GjUwVJyNlRPXM0GGciLUmCzCxLOBMfXdPgsqPsDgWlBRIMEd
qtvHMRpRyBo1bYf6U3b3vVj4DXJvYyL8eIoHOjHc36+1RO+8J+tYSKlAqIRxhBAuvTVM6M73rvZd
uIze8CgJy6IIZzInBoaal1Qccy9oOVoZOOvLywa9gHjuv7aQ3eRZCYNw9q+p+qBmGOaIqwl2gp2r
hxJjrD9OI2I47uFeMVkriK8HlRr0UEbD/SB6p/iLD6rbW+uzDSlouDxCqfafpPkvhRgtl7luTBkW
LfTa3hgnVBu6VchoqBqECGfKybdW2jBv8dVLu9r1591zwnQuRqCgMJ4aEwcUp/OOSkvxJP2hONg7
0wXJf1r/DXCF6bwb4yQPr71qJ0wOjKl0wpjsK2hRMSs8OuVp3MatIxT+ck8DMSUkohHoZ3E9OU6u
/QCwTh45MtCc5EMS12Z2aZMhTxKi+OGyaj3Spela6XwFz2RALy0aMctGKYAMKO5g9A0bt5P4Csat
YuMX84QL7e2oTSxxpiFKm90jaPwC7T4I/cyj6+G2RkBFPgAc1OsemhW437xDJRe9Oz7ScF3N4mYf
m6TrahTGDY4KwKqJmrfa1sMakSiQrGviM1l/JpEe4kM0FAQkBtOai+SsA3DZo4nGT76bGCyGCA78
tdgK73ZNc401dtAAFMnu1muq46RawYZdYLr484beSKtNyVWOqKOrBRP++YmL2b9mH6TPHOr9YfNR
VJc2h5ODfkLlM2Cs78aS+LjqR6sKNaE6WGf3G8xcEA4NBggpjqxSW3mgfp2TvzfMOMHTvDUbE43O
JixO/PKNNPdzPxrpLRkLAqKjswcBkrsh6v1SVlC6Mj5hycxjakVd5qUH+6niuq+puWIlTRevfCqu
THFKmOGSjglXCUVjk9UV59k2q4HyYOsrXrGX16QR2EwEPwM7Sdk4iqQUUW82P8MYKrptusWi/8+O
xVDeRyLoZOA05W6uLcnFGkqfSiRqkDuVkFgiRsOz+LN5tkZq3hoYQjgSJE7so4rtEj+nDq+/WYJD
lwFIQZKNMlg4zKzhHQKKRv7ZL2+c3Tc0Ft8NS0nTwqKuBSxNGM2WJIhji0A2bY1x9nh9/j8FxO9n
Ak1QlDXEMFKY+JEg4nUS3Knsd618oycyLN43Z06BttQg63fAFSyEKQq11RWBc97B7kORYJQ7AWK5
lGDZHMB/++3R/3UImX9mE4tmbCKGuwxyjA/wLTlljVZ+00c1/w+fIDwe6BSJpMcoBb5xLWHMCRtx
1Q097GPbMwIH4XpMxeVDMsUkCl+64AZfJqN7Sq7kRsFq2GrlPVC3k9SRyMSOVT1LNue5IYppHdRp
G6G1FYVYvCdOexuGHoofk0AKLp0Tz0Xwg9EvgSEfEuYILcRHEQjTHNi2MFtGR1V4bmpe1nXBLmsE
iJ2yuJBQwk9cgfcJouF67sMVwBFrZelG/hDz5/nnY9w5ZbELgu5GIHf7kAKzkJGtEDwa68fMWtf2
DLl76DV3jBaEWKx7FJsk0r+aZpIFMWHXimwaIHfvW8chD4Fi95jQLCTnMzP5nJ2qIWgPnooxuqCi
lfcgsk5NuZXpfprGm8F5CdukDjiQ89h6nQEeu7JKn4L39w3GvduNy+3hMvTsViqxZfAWjAswVKsh
HxAFAaGSsYsKIfeM9cHlF5vKUYoE/9cOmttB/2DLrtLfCxfMFrtmGy3KOM8eY/i6y+YbSQjVSQyv
l6AXg8zOWqrrKRG1CN3tVxQzxmwQY72MDHVEnMoNvY1csc3l1J8qtBIR4OX0DTKv4tvXLEyXgOnc
MYrDmF+C0rATbZIa9KnEdp3ct8v+Wf0HpZszlH46N3DEMU1eRxsIp8Hgmd6E+lNp9ioU1NXrf3cp
clB9vJzkzsamffYqS4en/YpBdX64lTxKPp6bWOmwXPVC7STYAlvnffvuVBdf31HUDtWw1K62OG3I
+M9wiqMRWv+HZEgIIXVJ6IrykueoqD4N4/WwkvpHLsqIXE8vux1OytDOStl7SDtshapqN5isxhfM
rydafZOYRLGlIPs8wFM5HLljqxTakFU9WhrmN6FCrfz8jIu7hYVKBd3GrzKq5hF0cJxi6gBxHD1s
moEh6rfwVUgRe0NYOaIvydjcFQ55uQ+xk07s+epZSxa9W060hI4T0qkayry6J8FR2EamUfo7j4qv
AJfrqJ8W6dWdG2wEdGJmzuY0q82RUD/rVhUSFhXxw5tkG50maTczLrHQE+1t2bNXoGLSSbqJmfhR
D1wsPbPkz4lQjE9ydvlXBEpJN5ZZ0TNK9+TBjxXr8QJc+NbsSYf4cP+OD4hT4GbdmgqITnrCKOZt
Njt4U4oAhllx2jkKb1xqI2X+ipYyeLwZrVqg85xgynD75pZfGgcXs3VqVB1ZvTDEzorIGFp8DbvF
hm1O8NryKLjlY89BwCVZT+Vc2kQ5gKpmT/BmhDwOP4aXmglP1/jLoleejOLInao40xUJBDfIuuE4
vuRWEAceDWhUdeWKZ/93liCd1C2nD1bBvWCLYg35QPfVq+bZ1TWn5NcKPYDRdE0xoqWmU0bURT5P
E3kd+q23Q2kHD3wSKwHCe96bqH0PRmWFvszGKrrAVFxMx79yIIaIDxArS8Hkozix4fxRhfvu0xb+
52YL5UjbmSaGfhvKqjwe5Uw0kEQVBYxIQOR4g/CQhV2NXBhGBCpHESpZu3scytsnOXGGaqa8H3q0
TTJsEohuEIei60fWr6yPbps+tqv5U/HMJbwNNQggbOF3FVfmC8/KVjGgbrwjR2lFZ8Oy6JX+K6NT
jLcwSSRrRi5wEdbv9JgSTmKIBq5/s9C5brBy262FkHQR2eywJxiExX61ZB29sib+yQAu8krI4d3n
J/r1NKVke32nCEMRAbw7FP929rUDt3w6td3yJkoqAYisisMBJ0gBpq7GExhb3PxJhIQc7amDiwHI
iwuqCBSJby/sInq+XkomiN+6TdJWRorlDh051+MjoEq/g+uKy/dFCX+YXwmzymJcpMtHony7LMsT
25eMX22p51iqESHp3JVkphjsdfYcEWswVtm8YYzqqaKEA2Ut/qy972qx3rolk+YrD2jlckXxyc96
lUjLIT8kqHlhLtOUdJ/aZ9jwcLtna+Tn9D8e7PM5dLv2bgssi22odd4f/JDaFCHpgVKmIv1ClxEG
elmpp+DMbGJp59DD4cmYO2ZLSyNYCKKWtss+qjlYy2ALUI0lDvOVjEibBLAL3iHlJ14xDllJU8BX
GRC9+5G35eBxN/yRYEB1koYnL/u/9QN+6dx9hjK6oIOF0O9LaRB2A68F1tZ/y/iLnDB89fBT+kSh
38ISt9YS+L4sHf7Dr+G8wkmeo7AbJastxxPqZW4gmv4ds4jxB73o/0DasbTOVzJDq3WsMXgnYXxq
NklgFpxo7b3JMCMZaQYsmWUy8EM97ep+Ob0qwhOsoEEAKhdxT3vDtJIPU8C8zqwdoN5SOoBeUxpB
KL/PL4kDG8ehItKwvrwG1xJImEOhV+NYHPIAtHwILxeki+mT7bR5n0mKfw6AMCkayuiveMXcP1nl
Y5bLlNquIqCcqoLjGyzqs9SAlPpglDn2c84A4aTmC8/sN2G263KrhYKhLJOXOh3/tdftTSz9c6C5
DWhn6XdmvJBASHVUNQCT96Sh6i8nfUGv53be3+WffNme8ZBgZt71hodDvohRi1Dpn8UPqi5Zla9D
EtRF6SG4QumXmxXbIV3BxbiH5/j1/kg0Te8ndDalTsYYHyOpLHgmHei3Td8lw0PqpWrOLeRoSgaL
iPpaTSleuR3GLsQTbZng1J+Z6PKcygA9RwUcjADffON3OlRN+gRWpV1mhQxala+vq/NUslPwwvNc
OxafQo1rzPQV8MezZ9kBt2Es+HyWyuupfs2N8baOrb5VaR6TDtGn8La6zLmIQDlQvGHzb3NPYQG7
FHqMWNtSoZgTg3HYd2tR8eCgAVgi32DS3e7hwGZThI+HE2YsPphM5AkdnkVQyp/UdyUQ6KltVldr
3UC+JaqW5YkvCAeFPrdXG4D2jgKHN9S1FCt23LFFIOZ5VfhSJlIk5WpxVjPNcnzxgVM5uUBoEVc+
q7PX3Br+zFrz3/6T1qH9c/FLYt99BSuVl7ju4uJwCov9mZoV6ANOOww/mFwk4L9TDUgbfKZVKrOl
vmK2d1fQhWDXaGnLJQSFbERQM2cu6AmtSy91HCTPSTw7QvyAdD/YP8alRe66vvgZkuDcqGl8MaGY
GQu8M1UdNe5YAb+g25fl0h/Z4xkrnxL6rwlo1bYljB3e2NdQm11Cgyrx0dyIJ0XYxIytAmMDtdbI
F32tlrn149UnrDA2ZuJNWskd36/ch6qLwIJrvPPioz+etDLkIgxDRagMvltCe/XhyUk7EgqJ+kjm
dq0zjIpzkCI5kbEXSI393NryZD1llBJ9b05bo7T25H4p7RlNjHoKaCZKNkv7xVwBd1R7AjQDLEjC
wvZWRmqcqNLK67o2ckbJW6pfPr8PHUfu0BCmB0vvTLW2zbRIuD1RVJtvWh0dZ2fFPPIqJ/PXP7WA
vs7xCQ82xJYAUH16Z1J0wy2/kqLqXDyCImr17e+oGP5LtUgmOR9RB5HI+oxx/0TYbABLn2hPHvmd
7AURbBvriW83wswL2grQIoOqs6XQ6zeVcCnBqXlxSGtGc/rdtPmSgaUL9MDvA0cekF2mNJWjeMq9
IAlVXpKwb+BjKlhjsxgHt8IF6wh8Ktbv3KyFxYEfKb371lKssZUUl6GXfjA4wIVsWtQ/m7XHBDB9
LiJbULDVZjNfXXeKZ6RqrNZqfnH2HV97jxXEISxTs2s7FpDdFjSv1rfWgPK6u8YLyeTQMk4VKqt8
d38TR7JSxYGJN61lFH2+YGfm9xIBoFYIMl1IfuEjkUULdbhzmIJjqGuRM0Xf2abTiKpneTo4qQAJ
C2IkdHWS5oq7XsWbW4lVceKfqTV7ax9ecjnQ+Bq4RpIQPV2T82qgAMivSuYDuKPwM8Rl1Be+9Q38
FU0aqD8uitoWg69pZs5nBYi92NvPJTv2D2J6WrvywKRVlHoaUBnteVuzBD1/AXkKzd7/WJbMKxqb
sjHyZbtjZ3aGeZ1deHmuDnS6vR73pDCwZ1Bol+1FEOzbekA2idBir0QnfEPgq4VnnpscdsO10vO6
alFUGcxVM/Bpaa+GKJXOQqRU1+CYesbfFVBjrGhNXAbWJgAVwKIShR6COHtP1tPaflxILLBFHj6d
mTLPzqqlsv8P7ti/cr1Au2Hbs6+D85jBsn+bpkN+8GbyamBmsWCW+vOArO8Af/Nr3L6uWfnR8Zlo
smAinajdwYPic2hHpM1MxXjt7hL5NAu1eVWVUXplOf/Hz8DBYoefwXNhRYXp3gTiITb4oHDBlFCi
qBBubnu++7pOG642/uYZ2BDatbb3QrQSQlk7YA0g3sTEaMarHfC+iVltiQ3OXCjk3kFrzezYoNIf
W8wdGPslf5pk9+yAzJjR0UbdkEuWYW0I+RhCjbdgikEjRyFdaHscpO5x3t/dnVlfs+C84YRtubwi
/TzA3njoA+W8vmAasFm9+e62h+8zNn1a59gNrcM78bU+Ij9KwPf4u8zsIWIurikeBtFQoVSx0TAN
cLWk4ZtHIFf3nPNkfZ/8KPJh7L9e1qJRoCRSjghswEJOKW4P0gwTB9UOPigcYhScS+CuyZaUyKAr
SmCBhoq8hEE9VTrqPtwZ5kIs4I7vU9UD/jDS1ArUHnbLEXxYybgOzF6ma5ZWjyx4C45Agw72+79A
SufHl0WINhsYamuLSPsyPIq+r0iPW2VzDFCoZmCvjbt7jcTEBTcF2ZRVD69/l5QjtPqLHIxe31CO
j8DbOU0K7G6mSNSdIb+9RhzoIWXwvpQlKgipvmFUqq/4+0t6NMTo2Jnis6qI+Oc/QDYjkJ5iKFUQ
87vTT3b9c4EhVOkR3GnYDpHAyqxblsOkkVA6jhRYtQfRpzmc6GxA87gJpJO/9TMGYA/AWwwlYVRH
JE3a1EIzLHyoLJ4ESjGz1tim+8NPgOSp8EWLw2JVKoXtaRDDyj+Jlx2BgwfRgDgnKF0Xr4fLZY7x
NCKX35IWTKQJc/QJADxviXiJqFaGDVqBrnI7k3LgO3T5s0yYeBCvtErpEZrTblG1X1iwD0gkgM4X
NijwfqmYLo+6HvA28Qj3sv90N5kjwstcfxaHKxJJ8W+BFVDnon5m7AcN/4yGhaC02sut8Fd/bTB6
FltGzmO4wqtqqlSvK5SabWNhZ3KYJe0QKXWoEvDnwHYacrzXx1zRYLuf0zFJX1sJDX/g/pBgo62t
BYhrgZ2yP8rsBBtvEFZbLcUAt9438GmB0XsKCkjzL1QMsbaAQaAmf0SGpk7TvkLhDOmLnf1icbUe
WEgZDlMSHzx6+H+hpPU2dECcVljQ9MqxPIZQbaX0FjtrU6tqWcB3RqAj3iULXbB1WF2nE/0oxI/p
PzjVgCs9NXhKy40ctWaLDCvG/9HnmJZiVW0GRPwvV99lN8MrACg3SKKIj9aWBk4QxJgBz7FLtMy4
ThkxT14EGoTVaFiNEQieA4idHplLwwJiSW48R3oBdXZQk6FnJecc8pnLObX50UUCV9Q8t77cY/a2
UhnW9oc8fM5tn6tBx8EnGTMSIUaXZ8XfGDRlvqgfH/WuftiMhEKPPUMknWN8MtnIVBsEg3nqwods
cxPw1UuvUr2pgZS93FIpm0zME4sT0gDJqquEjfoWt5nQiehYwNIZIWzyDrwIKyWPQQZGzFypoEuT
ZZL1OoI/ci/DhifuLQM5CxbULdvhxcg1qFieoTRbhHrXKAC2AswCReqRfMEc4AghLKASOTVYCVUO
2HM/d/fNJI29NXjK7SKp3k4S+q4Hl5AS6Mm96rIOq75BFYLFbUH0UpbS7Hi2DbUJihGxBGzu05k1
3H0VyXnFJkNbpH6KpIpZb8XXsIOhDa2MAzSa+1lPI7TsPwltptow/2Nv4wklIhyJffYgcOcP0fj7
bPAE74NZ9A7lyvi/8vWS0pE4FIOYQpNtZR5jMgXOq2lREzkpVLGDK8EGMkhppaMe75tOyD67Vnez
s+wntvBFxfDfX5ws7ROxJ6UQgB+qjm+h1hfgvEKgZthacShMrcgOngc2AJkKkfGHLJUB/RHvILb3
mnhPiCv4Z+vbFgizNw6S8zbSqkMEMhewRJyMPUkBG+8oZD17jbsrq5Mxdu4w27soqg97zRaGIKoN
GgGVheAe2koeNhITiUKtyryysKxjnoe0hK9ijLvEn55O8YeS7wcMtn1qffY165N/GW81XVlTOKZb
vhc7VIvf7rmGuAFebT665Et2SvRoLjngvfp85IqXJE97UlAQGppQwERPN0iL+1v27ly2SI8+ow5a
e9pM7kYl/1xo0J4+j5jKwgbm4CM5/OY05wdtoVlKZnJrks44lU6P5AV8YrrFk2FLkFQ+e8NyZ+h+
Ye6rt8Nqg+1171pxJw05P/r/z6QM4Uiy7Ov557fhuGuFg/efS7/tuOViv40JsnaU4Jg5hLVe8am6
ZrFFPuGG7o6UAzynqu/dqbaKxIFKliifkrBNxg62Ep83+09RVPy/B1Dn7laX63c4LEuCWstWL8Gp
3Z5brTTY2IBsEegzeUQjXrBMRc/0LCtrEyXJ8vKPlCdZEqpJEwYtSmRobpZMBZu2kvMMGKuB/kKG
HkpG5NEtrWq5l1WIIUFT4J0Vf/PWug40aDbfaB7LCEblTVJ9PVQof82E3dH8oX6fZbfaXX7ZL5tt
CsfLSS22gjRQ09a+LSljDU2W99HIkWuD44ATJQlcLALH4TPkiy+Eh2xPR7s3kJJyWsW/NsRhbzPR
QhmNZ0RfRx+iv1myXnqa3KqT46kAEDfBPuxNddvIBAVGE9rBxcifezs2MckcytPkrJrxGn1F+8p1
y2htvUBRpXKS/3xpm7yX1W1BY82zPBOQNcOd3HV6hy0RoxPTWh5WJknlGNiED4zuNRKaPblaMlTK
NJDt0ONitTJOHcFp9JOADnBsYQTySXpB1BXXI11xDofeLJMME8vfLEdAkNCQovKQtf5Z6gXsOAuz
7TTaLPfeN7vY39aaMqBoIWtAaJa/rXxXF8HYadXCTi0A7zH0F68oZ4/5hc/fL+WwQVPijcVtVpBd
2JvQq7lleuYFb5UYV9jytuNlWGZ74WCQ6GbtOEFSk1cgQl/TUxE/nfoy1uDetpZIdHW8uV2nq9HO
R4d+C4gGmABSj7Trky8ayd3mbjXRc1hE4xTAKY+TWLetMWKNpWOpnKm77fxoWUsTpdSYFFt2uQ3t
DCYrxU2MVNUP5Q0OU08BYfzqCuS2LdqztelsWNJJq1TN3kVg+JGZMOwdbzYpVpZOYOU9LjWRomov
8C4KazD/QQ1rloVCvo2SnCIvh8u+6Y6BiGx/JavyntnCHvPpuWt2Z7ewPagxtpI3CDfPls11WtOA
vYeY2UhUzgYlCK+nzZOBT/E4TefK2Ji9GJBMdSHgZm99rDniPcGMmxkFS47f2dsPl/i5fS+qeIXE
GNa8giYOH+x4gSa2Zu7x7iDG6IdNN8CqgGLacrpMZRdajMU6vX03yzL56qrobr/xbsXZIl0JF0Jt
3r5/ryrO2zfHC5fEKYhU7w0+juRcCNZWgO3a7tROKw5CHUWlpxdCmPCWEIlMvkHaV4a2tu4DwfGT
ASBZCgTQP417zbmWLAGUjbrPf9UmuJFP/252WCbcqBavqcea9hPPHKXyPjn9m7ocg4WYNm/pvocC
hnKUmC/RVlm5s1zdJnkhsBiBO6j3EFcOSu2V3pREQh36dIB/jmbJkXp5T1cIf471sFAtlU84MNr0
IJLtDcczjtLyjOTN+ntCHoxoFdc3MTios/lyr8wvP7qJCsr2pakzeuQMJ3kDPM/gJgOHKcoIuwVa
FFWj1IwCzIfBmMrm+jefqi3Zjul9mysR8d6kLp6BPcdOd/NDoe2z234MKpKplP9xbhaaYv/oqlv+
RKl25RevJeFs3ij0AqYMv7V3K6F5em2nFWvQldIXqrA7SYsh7Sp2lWXoBeU4qIJ6Abf9F2nM3M9j
KZtO7WhZGKB6zkVDopD0kvvPFlEL5WfK6tMOnSjWUUuRT0lyVPieyihGlXdDTgjL5HzK9SbNNKiM
3k3HjXxOgo/6c69xmPpnOaZmBqY0o0iXT/eT+TaIZZIsp9KZ4WH8pJVOGFVMOFVpO8p3NjS0uJzt
LPVlBun7fxARxLzcSHjIPPkkW7hyBMG9NWPrXEtiUSZxvw5TtT39REeq3uJr4+/e76N9qxRLuoR6
8Oynidn+p5ExzxmniQ1Qy7HnIoIw0IrTT9dtZfb8a+RwClPPm84ilmPfhM1KGEn3RcoWDa+CCmtU
t7weOs3bglWVbjFCL5vDApdQobEYDk1IQdniXWrqyfo9Mv1PbxMYpfr7nUGCgzx3UIc9D2J9tadg
2rnerhvy+jib+FWaDdFWTYs+siUHS3WJ22V8T2xOZYGHHnQaLUFPD12d0nJagbo6B3RjigZlcV9v
GX8+mofLCzZYtRj2d0yoJxzuaWmxB8h3tjLirNYeu60nLeFiQL8NJZMQTowvkyUbQhP/8W0wJ6Cb
NRX3xJ14KFdv2MZtUNFyqz6piIZ9H5UpW2+teDDSqDrhdx3eDRMR4ZWLkZiicEcNOHZevLQksioc
4vaBNcWePwxbuLJ+EksZHwGYZZRFL9OhZJR9eYyuzba8DLJfPBfjImg+KcUFgCK9gQwwTcx56Wnk
Y8cMjPuIhJ2s4r3GU/T/YHDCEobCwDUwZDQakjLCTdZ/gkzVrxKJ+Hg9fY16kxlp5vFlklFcBztA
Y6vMhyHBHl1ZQf0VCgClFwc07tQ+g32ydZMQhWUcdX6mGpl1rCAoUMOo9TSpnFYQWuOb1DChx837
j8ioih4o58HwV6JUuJx4JslnRkxDRpLLXVEmpA+eAI5j8Gc13fyMZWzRsaarE46Ou9A9bMG0Ae00
ahZ+FXDhTTq3aO1M2AaioETW45ZEokZDs2SoElUe9cwS9wVJ5Y0Cc4gWCTy//cooMfjs5U1wESgY
M3fWJl8Pbgq1R0AKS+11xNGxbXHCKIPX2C+c1lZjf/AbnrJjg9tBQ0d39sdeMiwMTB1maE6A0yTH
8Q9J/vUscS3e01wRhNsBwO9bcN+EMkKKtcw7jh5g8GrxidX4rJsXpyGon2S9VFkPvn2OvMLYfWX6
qJVs6Whsl7LcIqIM4OmD01ftgEOc7+C3emY8LPYqzwYaztzrCPxWnF1dJLy472MsiDYdGK4YY+Yg
+cgmSyQhe29+2UaGAPuQBOKkQ2WZKqGZ4CvJAooad+Zf5Wwwjez0BiCQ+P6VjGDjQqGDdXnyTesC
CL9Wn44Pcd7gHQpq24ejjUJIPKZ8mL64FFaZi5G2qwEvU560cBFPGUdD0sRVzeupune1ccMfojtC
4WQcpnRRtYoirO7UWxMkSqkMiCsB6Op5lQAgH03aWVCo6QkRhV+I9jqQzyeZcEHdkBXmVkMCrgiA
hX36q98tD1+Gv39NJNxiV4SfdJkwovvSHXjK+ntYk3UNHYEGITZrh6etHsKEsyQ6cv/GDm302wMr
M/PXpbSwJJhOg1kyOW6v/GR24FN7yPrvA5jGBhRlNv23iHoBBo578mIdfNPFdZYEPNSc1hDEMpIl
4XlSoRIOtBkeVaQgyf+/bWeqlNAVQiegzZKilnKhuB+RxU13ei5UArYR2DrbowKzx60S0+6/BiFY
2MUNQlcQJ1WbOFIbOqLshJJTlMp4DGZV5EelWk9kHX0usg68GHVulBj9XbqA0IUE5XKqwHhzZR5f
Nn8ThMTrP0rwdSODvmenxUE204Z02P0aXPuUVj95HLS5eEZX0wdkNd31rA8RJUlIPyKu4DjLEg4t
gWrxz80h+tN2qelPjxOjLHY1/MI6lwVzGwm3sIVywu+HWMv20v6+VPyr74K2M8dZboUhRqVcOad6
By3xFo0kJgC6N8yCAnpPCRxXxCIsESCTZfvYhOysF+iSN1M2b3vvNr9ttiTyoY8GgrT45ADjkvDe
G6f7n4QH0BDv2LHxtOMiUCCWUxrbA8JBiWwbrP9PGkLXCfZUbWyG8C/E96mSwSL7KVsBaIooLhj/
7KYa5Qo8sgj6UFJRa6DSOZtf1Ey3jDIYWg4DZ8uABeqik+xrI4idF86xoAuBC990XAs5ft6MGkIa
KK5k3BqVTHXHj9K19BSoIUgJFS/KjCXAscwchzzT0E5/JUKI8IdadQsiTf/e3B/0WPyMKsa1G7qT
eQBdszVkrta44wP70Tvd1hDXUfWZ7yyxhuIfi3chZdEyiTIDksot/MAo7IzdxZhB5HDGuQld9y3l
HFxK4dUJ8uRgme93Ft9ISmKm1I08WLdlx5BccxiPlxQx66EphbCjnvRF+zYabuH2KabqEKtT5KwV
nLL33TDuhHSlzXZEIrsPUMDLM01HvzlrKQbU6Jdyl/+ZcFJLE3UFHe8fDcA2umAub9DTtcv19Azg
NZznNInCEytFdnld1qA/Hq9u55CbgtZpqVp2KEHJ3iDb5hM4DcF3FKpF/ZYXMjcJhk2c+TUi4DQ9
jQJerRYFFwFscioG4Pgmq1gzOKmR06bNuEBrw3OzlIcyaKKtAC7SO7vlflzDDfqG0uOv5LteBOpL
/nkJ19y010KRpJF3gSmeqPS+v4zH9CqIQVGvFxje5ARcHK4eH60H6nnFKDnVzJC5W7U3Zy23JKGF
V67/GTrPyxrFGB9FKQ+QAL0Rfe2hZVzy2Jz9DyWzeZdU3BI+AgB/RcAWcmfLAVBOiprXAKx1u6Vi
prehZIfGxaOoYJ1Vt5a9c7SqIzWH1uS7RALAm3CqRZ8ypf5rEzRTi6DndArWvgU3hCvDffs1FFtO
TnkM/zCw1MKrLOnVgXAUnEBnmRudtoIcU8ADfRXscyhZMy5lHu+Io5srdjjQ4gcxHbRlZMDqHiPd
CdxLkVGZSCCnGICS9rHn8vr4TLUDFmtL2fMtMkQ7ym3OvB3iibAqlD4qvnrjk507DwqVHF2kSnSL
fxXm4Lm1DawMRG/T74w+bVyovtsZ2idgZMg52Z5gd+JE+0fnBSIUgiAzOL4lxt8vHwC7dWmaGeDY
15olmlk46tG6bq7Md+amLz4gyWU20pUQ8WCQe0kNz7U85ZBq3ENQFkfLjt+ZCQWZKRFez3MiBRfg
ppopJ8eNCdbFKhltvb4QxiR8liwQtEkNirEGfJpDFk/XZYZguA9xg4x0uY1ez+i3uS9i6CTvr6DP
K+1pfMdSEVuWZa1IIUQdcRmVrkDGi4hgnrhtWcK1Z9Rtz2aLCGY/GVZVnNcgQkTLpXXZG8GQ9nzW
1sd+hbFzaRF7iCxXfo/y6HKIO0pNT6iRi9Xv7iX83WU2IrsiElJ0K/5fYTe2tf/HB9/MCwUiGIrk
9KZs1KiIUmKH6zoSE7YkjlNerwONGQZ0K+0O//7P3crmswsR1El52pNnyTpL/gLJlYA2CjinZAQz
3jvbcifq3FWENcNwOmDDySkDhl/4HLa2KxLj8p6d9QQQOJiWuOyk5PTA5kfV7AdDE3a7Scc0uvWd
3HKTTRUxzg5Niz1lc+c7a5wEsvv33GGnVlTBDUG9nD1cKJxxZBjXvSDTg351gHECdwCYK2xJFHUP
z+DBuP92q0TDkR5RuXjrDaDbMq3+DyPHgqR4Ie2ea0vl612VKBAJsV2W8MkSoz9i7o7nvJP+XmGm
zrUEf0D3znCAb7aD2WBr8k9ZRdlAZM5zPDADAlf952dZSBfOevz9jsJkODcO+DywaywxQinqmrWl
MBtK2EUNSwzGeaWdqyzfXEmA14YzyMFN4oMeZzDftQKjLnR3WZmr/KE4LG4NNioTRqLvNK+06/AP
YizTmA+FqYiPb/Aos3DlxxLnnNbouFXUddNZhUPTG0H9y/6C8D9Kxp4SFe8TbiAV+jsFA2Q+8WbL
smsrjTj+y/NUViW+EZJ71NiWWt+lLfgA4E7nzAO6bfb9rD3lFC2GhEPzklLR/UQO+wMAPowDoA/1
9eQu5wemM1SVvluuQaIKByYim+82sU7CDwY+NErzioTKi09MGRd1lzko3uBk0N9jKt/iAyWZBMmy
W7akQ3VHyleK1u/41Ul/rbIqzwYoNcQPGhEl7VqSHKYe491C8wTC0zJUr0oODz0tX0J4UQNmV7Pw
UeKq7cZDWsezrsY7Qcx83zV0AZdDr1QhJdzDoFEcNBsl+BvnND7rS+DVr1noZo3NeFqwgekgCwgB
P8j24uA9hZ/L1esPxJsbvWjVsePfXrZnl1MWTuJeKcu4+tocW7BLUVyQAu0cDP6K0D6T451lo98p
1JUpJHuue8D1vSVdwhlX13Lsz3JHY/gWo1kh62nrHYfCHwLz+oOTZszmdcF6GiAB+/RVg1Ks0q/v
yHe34b0MV6Wm2lQJAESK3/+rdUk2pb1Ux7VGfFBZ6EvQ3l/j0vmqcDubL81jz9O48YFSrT8eTpzJ
eci3FuEBRLQnwWhguTSp0OKQBKYcrS2BdVQgZ7BDUEEU+KzK+03WF7SvvrvVAHFYU69OQRvY3Wuq
IgODBBtrhgF/GwWYLLMSy2vFABhizSf7NVCtg7H1GN63HMbdtbu5CRXW8E3Bk/dyj3sunH3s1I9o
A1Qho0QDWokwEajcGMCcdUINtPsqlSMquHrPHjnWfZxO4G12+R2EETBK8jrQ9Gzzl+Skp4PIHq/L
ObXDv7EZkXPgoGIndhZi7XngMMONGzF/W9LP9KzgmugolYhqzJXp6avTkYBy6DDlJNhNWyjseMN6
liN+VzluVH3Fa2QRqCHD8PiX33Qzq87MbggakKqcGkWMMEVPuEqSqZd6+po0MlED1xkiL6VGWkVs
+3MCp5kI/8aAJa90z3lomxfto5mllcGtqxFm7dXHRDA7X3QhELAt2SJdSlF/0n7G054J8bvlqD4E
m/UY2wqU5ivMekobqIZuiOh4bh0GLH2VCMX1aho1g7iHpolDrNhJI+ecuFIp5N/PuBQ6InR63iL+
9R5xsKskaGajWPlgQvLs77RtMkzUbIyueRtPZrGe2nYvRYb+kgHWQHEW6bIdjnhhmutXOLYcMoA5
dgeSsPpfsU0Aw788NtRw5Yx5fXH9qSabIkdXr80k17Y0rIWhoan091aX/rq0UyvqAB/zkq6oy9Yh
2kCEJD4+wEUtdOK/rPmJdLcJpS3I1LBhm+qgEFsPCDDAkNMxr6N7GOVS+MsEDN0pZmPBP1j7nN3q
KXsQlpRwRvpbWzwB3hoZ6NA5iY1rq2/tY8X3noNfz+1fD8Oplu/nEyrg+yvBCHW3/SVzD15MHx3F
x1relB33nD2MR/z0NMDYPAbFRq3mf/OBhy64QNS72QJjuaKwhqy20MLNwZlLMzsxtmoDmsP8Op2I
kZfGxNz1SZfagj7rFikJt87A4Lh1JFGu8CSv7Na2sf7BPiAWU7Kgobg0UznxTkX9OpdGxc5iP0+f
Po0qEHx3X4Hlt1eoj9nGzLvkQccMTW4vgAlJxgOjtEgJSpm+ze3GkfP6gK/8xND237e+Z1idEi2M
xxz+IXw0CE0AN6uSUrPWac1ALSSYWCm+rG6JpOywXiOUQZNbX6CgvBX+u+kRsLAclKdY09kcTOB1
+jOhnBb5rzFN3bivG2VuEr4ZUxSY9z6ezbgZWKU80xOcedi6yD+Scw2cdsJzkn9YGO3SDvJOJnjv
7aNIuSDvKoS/gKcq/teBnZKRfFKDvnumZCLMsR4JbWD7IcsZH/O+t18VrHwY5QPv0QgAYd8vN2Zi
2NL8OlLvd3xJZD3SlR6LmY2GnrB8HFKJyMT3hhP2pktPum8nB1oT+uiayOy7xczFVzJoDZYaw3Ct
hGqCdzBjox0wz7YjPKVB9eDqyYNODrctGBnz/gqBT+MQIM9z1wBOO6n0fRetFSlk/PdnbPDV6Pqj
vM3Ku3gYnNwifS/DFLVIp/y24qN2UnVCz7RYMstB/6x8gozdm3NbQKMWoMx2+I8VuWsektCF9WQ1
NT1LCJPH42xgeviE2KRS1BVO3n0lxcry2rerzVqGkpa4uJg+HJEOAfHT+M3tGUJxrLA57coL+P3p
YUgojRYaPEp4o8D00pq/Eh8sR95Bm9r3eaDrXucQ0r0EclJGxinZD/qe1p6/JlYdvG+1auor/vZf
uaHsqzEmHw+eU63DHlaO7uroUlN88gTDexDfU/bf3GDc356ACevEP+iTPlPuzjID4H5CgAriNfaM
BmQtsV1jHuSUNvqRU2zWxBEcCwvMHtmNP7WZc9J72L2uSoK7y6toI7mCBPCWn3x8bL/sq3qEMD6d
Mm6KcJMjJMJdIx88H/SyvHFM/LnXYPE+J0IToLss328L3gdIpoMhh8jsG+xLcYi2M9PDaCSbGk4X
WGXHGUFqyUvPAKSe36w6ACtjmBegZU45Rqmf6Fh171O0tNQHRo/cT/Up5ZxyYRWn9pU3/ODbPILR
Ughket/GO2Is3oBGK3avJd8wGnyF+ty17FeEnaIBm0w9R5EmTkmxgbCjMyFQJ5JUuq/U/DgVSves
ljIEa2YtABi7k3NSYS/zf7KnNDn975nftCqEEKQ8y+tLizVnhTbe0+WHLIOng0+IsEpcELLInGYf
xWXLPDKsP0Qk/XSVcvTzYsHSLhcCOCIRdTkb/m0OSfJPVU7heXHqxNXjycoqMwwCR0SZ8ck1oCXa
8MWQpy01Tcf2ksLi9Yl5lsBR5Hua3SyeXLhCZ0B4OFytQojJ/i2GQ5eMzTSIOLvtSicx9acMsuz+
dWPXTJfeW9ZU5MyaJ8XydQwp61x+kOQfcK7McCBrw9oI3V8Djo9iCKoUOql3BsDORlqZdtC6kaRi
FBE+oYnnghgbWZIpPpULlnht/PzdpcsHG99NNZgR2Pv9f9ZZ1On0eMgHvP9jklfHtFSeL3W8noME
kwM5EmSbtx31AVO/PJZHkZeLLmPGm4A1Cl213WA6JOlVZPJvLFHsBjeuLQOGRNsvuUzpl/CFHDtK
532R8rYLnH/UZ0Be3kahfIDMYU58ALcYkCQUTMPGqSOYyAO3qRa0PjBH0R2Ci4/k3lsih+XqpZMV
bqIE1IdaR7czSXtAw9PH3Gd86GVQgqUwCcfH4jeJgja3jk2vTtT+us1oQ2qYAUDDwJ5a7ICNKENQ
/9OHQ08OitbdLsJpp/6m3B8FcIiw6cENSG7qfIKgJkG9fwSnFtZ3naun3B6kXyKA2WqZt9QLsZAi
VJffbr6Bsyik/1zNcDZjZ61QOATxcYuN8+8LomfmRQgvfT9TEjljegqewMzcQ11a7lKAT9qtU5oC
FbzQTg9trI7ndMJ3qSXkmlmQDSLlasmLKm79+S4Ka7PpyZ9iNdZNyS01a9MLoqLv/NHmNARSJWl7
w64uoxZsDXrD0CKgcTPJ6bbCM3psbnFT+GK/VX9gTEpCOJSiWSZvKQHyR7b5V2ECc5Y4CXeL5ehA
ZZmtX4CkNpdSdjA65dXAl+gxohuu+pWMVeVrnrkmElSJpLh9Zr+4CpebSWgj73MTNfjPSlm7zPw8
dfU1X9qcwes0XdleF4S1HygDLgS0lW5gI7YOZI5xohKSQS2u/RHeYZJ3rtCCzGxpt0sCv+u8NcGY
70Wp53PfF6WW2rur4H193Kqc6YbX6i4OoClbHlPNv/RYWfbmplfomYRB/412765p2byFMj+yImxO
4tK5yF2rIcp1haz/nMD+WeZiZGpUsRndJDHa6PwycozUNNS71RowM2kC3LtRTeO2q89R50UUfbo/
dr1A2SMalB/8N77FMcah09JpOl3UeYFYLOEj7diCSq7/vAYAlIQehPNhYxoyYwQ5B/w/13vurV/r
bg8Bz2iB3aQ2Gn+rshXNNktzdNITLfx4JiBgWcARQzqhlq0Q94M7aLlgX9IW8VhewtTyRukKIqeA
OBFXj4W3o9QvaIkes3ArajYAoJ/Ts/Jf4/ygeBEwVy3rAKRpOUc31EDjfwoK9bLUPCrjoBczC4EB
8gY2DMuiRR6w+3FML02RIuWY1VMvEwnIndeqRcLzth++hczy6xB08ldU6FidDgvJm+jS61FQrjSE
9MdnCnmtgJcKbhhyUm4BGpEm8ctMudVOHHFzmYUC3yniALwLqlMhVJoKwXOt91p4HdQ56LBxq3kz
X7lWInra0Lkw4c1TFBpmkBFpaSP+z6lzkAWdCsZJmbhQCE2Tpv9/pwhC2YmCbF/LlkvzkRklZW5X
Td9BaBmL4d2aoYpB3V6I4tZzGIqSZhpFlvWJE9+8Yu5x+yQZEIkrhBXGjdxxM0BULoyhb7mCPeDr
QCzRCuabsGh+g4b3Oro1yaQjUA3Vw4SvQkm5XTEBpRh5cGO5prVqC4WVdo3KKNnpsO1h+5XuQOL0
yGicBji/sw/z5OtlxisURBt57N2Qs2g0jiSv4ViO7ZuQK2Sxkz6fszCdRFUd9q04Mk94E1meA96I
9XDxo08PnlOWrpO9p2tpFz+ChkVtjnQJ4kDuUNZW5o368mI14PnejtsxewYw2L2/0/yOW1C3no8X
iGNhljWP8N+e82yadD/g3x3NUqWIOZXfeTQcQK8NY6H76yoXAgUrin6DXHZ1Xpp9FxeFawvmz+pk
0BjDu1txDWxjULP4qqbfju44Rk6DKYhWBhdnk8BXnxhqTq4KEsdcdygElcGPz6b5r4JJDqCIWXHJ
aykp/xLVxyipsbendDfBb312kq0BkZ7pWu4923HKqtu3tgHNGT488lxwJbBsDWJWl1WHvHXgmmac
ar98pZN6qBAu6jLeA3pJSfVvHfsq8dqqH34YZiE2afMv5Mi0My7Q1rvr62EU9tbyT4SoW97pBGkX
kBwt8Muaq3uzMPbShbB7L3ZQ2vxhh2Rcm9N0QPmsBHZ8YT1UqLG3MXCKQuy/ZlzIfPEHI0eR6anf
l1YXIa3DCahYo3KdCXmFh/m+hrE/KiT2tFzaTzv9thBoAM+/SB44B/02D9g6Tl7wO2NoLcQk/a4t
Gp5Tl+rylemDA3dQ0XwSMIiZJd1xFALxlN1DvPUjKG5MYXj5L23A5MX+m0GX1O5Eti12FhcCBFwr
wHUR3ebT/BllJFcmxfIOTNaJ/JMrG35C2nVtS/ueFd7or60HPI04Vy1jszA7RhSUaGnVN0ki86qz
a6DBqf5i7BaND00iJKhJDntoO1czH0ZumE3Dlj/IYfRHibGrJ9CHBnnY49ohzIIgC+2AicS6i0df
cH5CwgzBumdSmvkrykODak5d+m56t+e2HGZ1U5u4J+Y5Mn6TlUCftJs1fz9Axsb64w7SFGVlriMX
emGkeYKoiyS79egk4U7isZhF+FTirY7j0RQWp+5GtI2VLGRaexuvAeTV9O18aA8+9kB6xuMQj63H
2BSaW25uaSj2HCl8mwltDG9wRkYOPik7DyODdo+0gwe5bltLVXvUura1Ha671hqKKuWOCP0yQhiC
G56xpxcBxeaJuZLxRp56wM3d36jiWeeXnHPfAZI+GHZktz8NvVdorXJq4ECRdrYy3Z9EvSCbKe64
NXr/Cv9xYu1q0XGzK3xG1bSVA+zemySDLwNY0zO5ewcKM+eX2Rf7o5NV13eOjBn5tuHWKx3MHeZw
qYWjjCL98dR+sYrwYTt2BGgJskSr3AqSCtrkWdK8krNPPowhMY8reEXaLyFVJ0Jnq25B10c2X7uc
H+yXoIWX4jIoOCFDgoNkNzrk1yIl8Jmpcl2ZxRATN7Fdze2DQ0yRn0A87z/gvTKa1riO6p3WlheC
w6U2cDaH/lakyGQSsaugz6BtNvt8klUbti+OZ431x4+Or7BBhlNDAtKoUu/Lbv8m8P265ehZWFRP
QPzd5b+TmCbOTv3DtzDXUB6cIoaX426lHBuy9XwAeksxyGq2Kux6sl4CPaIzYoWmlZo05y7J0xDO
crqLTOtaN2ohpwv6iEqy85/SbyEW8CrI4rg8jKisPP4wLExGr6v7bvz9fC+VAn8UDlsNO0XyBCeR
tATM41Dg9wyZErco2Fh/G2PjT+W7EGsNUu/qfMKDvtdwB6qZpohq7Ujnfk5gjq/fiEXGv7qdZvhj
cRflFo0rqi26PwA7JHw1Myze/StrINa6k/xahOzmLARV0mIUqmO6VgdgBhX+GDOPHqCivNCEZ4Qz
8yAI4eNji9ObgFj1h19RDbbfXjeHjVvcBkdFTN5YYut8wN49XPrgXR38Djdlr4VRvIVMCyWrJZXq
n/JHIUxXEKxNtLxkaDpX9/5zCvH8hOwTg0PC5RjboiD38uiQPm29uXSeMti1a+KnHNd0WWTA4pdD
kxKdLHvsOsQn1MKoqQMlO0IHMYO7xh00fY0lulrWLYBEld2ONSojK1/9gNzwNyBvb7Z++e7aqq0m
ho0M41b6DzjSYXpY5doPEIafYqZTVkwEgtcqgxGwwyHgx06Iyu8c+QQLoSgCM8raaYMNWSFdb0fI
sDn7Qrc4mYZPQAm9WbS0mxRJft7SuqDHSWXuRBqO+2Y9X2FpKW6gPhAzBPj+CyBQ5u/lFGFbn3id
ZFJ9E+PGmIcCW/DH2pJdkdPC7RL1MrmDGKZU32C0lU37JxULmcKolQ8Hhzyzn0fy914Q8u7tAIMH
UP1jTQNVhiCpOcTcYvHpBDC0KhJeRjFxamczJDKD5NXDPwYtlala1KjgRZ0jVcqzYpGwgPQ3WsxF
RsWU7RkQSHqtSh26oQcnKREmgjU8dNeyR3RAPRUPw85ir+tG+C7YHpCshnY/epKfTGgnEuWnqiV5
paGlWz/16saHW2MMCGdtpnb6sDBVa1bH4vo8GJovfRgGgxvaLbq+6VUwtADoBji/j6V8zazeBKU1
m6gdPGRcnZuHlZtevok+sgwtERSlpyBaXr3/QELICbWyHNniZdBsrYbCxIpWfREQIf745hTtgGtk
5MRnNyGGKqwkndoh/ATJ0fSkJF6SY+VPn118NguBurdhwllFXYIAcf3cmimvCAM9oPJLDJdSfwAM
2Pt7bKEeWDqrEp2n2dl+T3Q8STpUSudhnI+2FtNUIFpEumLIBX4EpHq6i4Cxmnzgbjcm+Ovdz6TK
qiP5Qaj0MW/13lMMJU7LV5N7jTMRTHc05iTgnSC8XRH285HVigGqm2j6MI8/vLS4t6HDBARopvfv
tUAhUMlUHPmavSwLVE1twxL5U5Qu6P+mR9yONgTExjGlcWvIOUVj9D2/p/ORgPps91/PA6eW2PB3
4ttXLBrmugvgYxatLBi5P2lufYLth5PyhFiG5lnuD6U/HJoNZuw3EVJ5/wTFRM8fWyH3T4BjbuI+
l1D8BmGU73qYBEOTC8f94rargyanhD1jjOMEUQsuL3bC0bNWaSfg8Pb4nOjxlwx/lbfF2bOlqhhC
D6SRtB1ufQgZlET3bt3wkNAEROOz3S5S4Hg2+ir2C9nouM9zZ4m22IKzDJmNtl+Y1Ys2Ld16VWKp
fLjLejCWO3iQwu2Aua6aBEQMnHewVVedigzFZRvGrPOpGMzeq273prWp1PRQbosQy52OBtaw+iUR
nlDj/ZlsfDJ1LvEbHAyJAy0b3KgOXXlCHO3lpdA0/zrVXAr3ku8FudNSOy0TdUWe+21Mo+Y64RSQ
nfGF/sqiYxmSDFwqwYByuYdYt7Ujh2NuoRpAuFqpT6hwtM7x1Q66avYyGJp+qiCz/2IsRR2XTQca
ZiUIyWltkcj9LLV2+aWX533v07Sv253w66Yv+CNGxBVHbzX7q68ZMVCA7CpdNIVJtnySkn8ueB+t
96xIiPkB1WCD49m+oG1jFI12nF2mRNvXUapKYjd+5mgaEUSU4bx2kX462zPgJkR2bB1LLZfmu097
VUqxsoBpMoLgaH5SCisQeUcc8Y6OhS92WC8MAf1RcB87OvmVJvM0GDE0WI0DFcuWgPPBhVI3wmpD
+KKukGcp92wKLFwZV5WWDc4EwoqbIGmKv0njxYMRWAedOW9r6U9r3CtkF1Qw70QTOPD3wUz9F5X7
PEk4EuLq/xErV4sOt6e38InVPcNlXqTgsW8mRwpMtFpIVK22qyCN3gY0cVx2fLWPdIEcAyARhP8s
MH/2oPwvXB6VbBic1ezYfnAlXFXOXm5KyMqE3GM2jS+rDpPtF7MmcD6cQ8w46p81Kw+/xjj65gd7
oWOOL0J6CSaY/nM+u0kanByuup5xhVlESsOedxapLlEMjDrvcy98U1MbmnzfUtq36ADAlAYMcPWU
W+uZ5Yyk9hbQqAnh0myNQkU7lcnNRPCfmkVBkDI0mdliGi+Xh6iUFL1MjB0FaLH/aFVZj9waMHpb
hSALcbyHkxXkA2YjT113XigN4V24nkVxs2dBkNh1e0Kc+nUyqr0WXFTipd9RFTtAEIC43UUCxTfC
1xTrhxvIpIAjIpwiSlqFVAQHBspVJC6MFXyP5jb8JkwNSIMiqnxQDLJqnVPMTI3TMWKvJ3o+1BEi
TzZjbsakbecobmZaJgCd5G6XKUq/a3UX+1uvX5MnRGt3MBv9SiUk2VZOZv3tyYrSdBmi/z9/eZUl
a6MDEFDO73DPHluli2q5vC8Ya4RGHZtWeENPgQxScVWPtcT/ukrsXK4PrsuiUj7MYRSpX5jxLfCL
FMeD1/vYPnr9ADFRIS7EwN21wbZu54dDMQvhsa+4kgNkBGQhSvpMBjQeRlk8MxC0EmMPMmF8j73v
yA7qT6GdG5WHURU7fK7WGwwJWfqvjOp5RRBfxJHjXlnkXpDyT7pkM8AplfyNorqlxCgs2zqyA553
im6W4FFevREoB/spBEZJwzZYS9AgUHMifw/LkhEKpauKyabLauwKuBrpYCec82RJQ0uTIFRbl1ek
2AUA763qYZvbI9QmF5XsldROR5O2F6Olykbk0DZc1qQ+4/811vgHceHzThhsReWh2Tzw54FdIudK
dtUAwSK5go5j0LLX/FMYvAowyy7NO/Tsttnb81zgRCkC4hWz7BP66TvvFlVlzuPaFUCSplkYstLi
kHhddDQkLVC+BKzntMPkusWCgyfUP4X3/V230+C8wq4QxJkOd9hjpPqHQ5bNdIVbZP89LeJlI0l9
rZs+nnU8bvWTD4KDXeZQtipng/4iHCcHqbA6VCnvkt0AVF39aGhSscQuFqMqqjaBu3XddfFfbslJ
zJ2kBcix8+ECT+CDWCNvtxW6kRThw8A4Ev/mrb52va9JBWMMLE3rQBqAGVCuEY95xW/F8lLvSDWF
sGlbLTT1eh1svQ5Mu55iPY54+7mqz9OFvQdwAR2Ldufaiof3WzwmZBFnNugxIH51d3p9DhA7xdcm
qcosuP9VTYkLZaaFhgXMgQf/GEaBDVEqp2ODLyvaHvz9AOAULoKVLvJk99jLIgTv+h0RFBWheZV/
uAXz0ABwjNZy3DjZ3FiTNF3p4re4OuavKgL0HRaMS4MSjk2tR72bI33yV1MiRD551sxg1v4Wi4gN
aaJj0xKsXFMmJILzOUcLZzXdOCW1rm2XBXjhdpgBSHTE0pqVMzgzlpgvLoFgzGW3E9piKk403HBY
sp1mEWClKk7iuyMYbycQbGOTP7ALtXoeOrKVw9iibhIBB6jx4bOFsPHc3bIQMpa1MdWSxpwlpGky
0WIc6On5SSNb0A2W/rR5o2YK2Ggam0d8nW/DDz8iZ/NiAvmrKd4wSRd0QP2pZs7ULgyBhuy3uTLP
e9+1uT27hMJzufUTrxmFmYFb8/ZvA/C+7wS4zP6pQVH7p3pat5Q+fB1DkANPw6+NRVFCEHH4KjXd
Ixc0nFUwNsvSnzj1eVteJYi/qMau7HWH8vSJscTW2VcAVGMSD1uQQ7025kUZIViN/vguoHpoHRjQ
TPqwrdJmmcKHiTw8CNjR9p9fl+ZV8Wb4BkR09wRe8h5nM31ohKgW2Nh50NVUFesJuBjVI4A0uS7w
MQMtaPh65wg/8GXBUx25LH3yozRGz5FYJzmsB/6VgBp5pEEDrEZm7caQSxzt3sCWaTgGLeLWLMNU
6O7c+0E1tg20+V5FKFahy9DW0aMwKiTbS6jVe9VntcXT2nR9nmwK1FypszsRk6aBeXXVcuywC9Iq
1xOlqddRtq2v4ul88KV3O6VHIVvLbbyQHSaokwpJjra/18u17KH28Kf3sXq57/95+QzHvb/K4gjl
JqenUv4wi6GJNO1aWf36ekcRBsEe57kqyjEjaUx3XmOWwQo+EhVuTeoU1hwafGxVY4CAjD2vUSWN
TyrbPDDku76JMJxXd7fXQGXoTFR1xuzriuP+8D83J8zCAGh3QcFXFC1zwsi3AML03Lb/1zaD3B8O
M72LRjjr9J43jJKvZbkFBIUyLrijRoqOoBCO6S+9pe2IMDIeI/5N+R24IPUhvaVSlaIogt/hUkY8
+IHgz2IjBcnenVmGrnyCOI4TSCIXZIig4CkKHDatKVVDVl1Z7LX9br9EnzM50bxXmkwVg08vUCY/
uJDLGnXp0148rqpPCngOphOYkCGve7OrmEYnV3qnHHnBtku/AXEe1p0Q1b4XhU3KHynlbS7WnmgT
xLIAU7yP5BBOL2/x1AN/QlfON7EGG0WyulSRYtcWuB3VN0bYJngNq4BOMyaYTT8DesraoWhsWCbp
uZha4lto/u5xbkoH/hPnVHha9HeNCdCqwhzqcc7WatSCSKktJPRm7IwoVsZq+GlK3OeY5XD3EiDo
lDixByhn9MnC5CkT5swdAjOKrkbY5moEeVU3Ddja4Rbf6M7AjrwfjM/JnKYQXgklS1GjyxyIGCiR
EhfenBGuDR6VezH0b1Fm0+BRm0lmCgEaWhNoyh9Z7c0EjGLyJVhICYXjix1xCpBFOac+ZNeOv4ff
FVVMR0AsXeBgerpPjL1jCJv351Vl61o+WKU1UB38gOrCDufAqlTnHJ6e7fTBI/2kICUyCcZbgyDx
i+9qpyCbATbp5dFjr3Ak79tstYFYD6tawfnyGRK2id3ufXdkrkwhl0W9xSiMidhglTMKQygJdCig
Ug6jFuRHcZCzFSqJI9RVpKow+X628SJVyQPmNW2t42Pl/UCuVC+2tGZ520TH/8t0ExOjBMA1X3pz
MUaB6t+HPIlwl1hlKJCTh3wEiSk74WDQ/zZRuhIQWoZwQrdB/QyiFO5jgpgfBEhqXpfh2MLZ+XPi
DonG5BDwtNb4oLIyaHE68fqgZ/ITpknhMGKgvLptzwJ+Y34hhHz3H7lCPvGDGgBzkG757oorEX4u
+QCe2UV36xczvB5jR5uiz4dsiqjmAp4xkK4LZ4qJgSfSiQqNWBTyC7Dqvs8sRjOMoKljQcuj8JbU
H0et424dhBYGymH72aR8gjWo6pdUa/xk+YcWpXQl2mW2gtGZBmk1fe0GWVPh/syWRw/67ydnWT2M
iyFoGOymrbxG+dD5hm9pFkpHZwqT2SELi4N1zGVfrD3uWsp8UqJaNZ5TiVhSzPKuAz6W9FXgMKS3
8h+NOsupxcAOQb8rV/yryVvUOa59pfC54Sr73CRk9aVOzS5WtPd4aFmOc0yPLM3H9POE0YZvIIFB
/Hhg53Hbre2Wuseea7adgTusoWI2wjt3mZZqTxrAwxKxK7/11L09f/zMejcAxDY9RlP0wRItjQPR
xicNb6jaNhJSTzJaViUcBX7plSGaJAUnmtnO6Fk5I8shlVjvWiKOt22iRc++ke3WjodvwAcy017W
SJqVrEjtrXLkiMgwogixmmZ7xXhEngNoGVsKttzrd5qEvqd+7PhL2mcCSyq9xDHu25Efr8USboQi
hzuAI3I6/Fwb0FiwtGfOkQlt0xD+oQBQmHYHVOnW0vZ5yI5Zaq606fPYEQLFyWHBLoI9RDPKX8Py
KFEtBrANkARFTB1Ch7gJURHK1yTqjQfZOMkJFNQfzoXfg1yXpXRtQl5OnFnyytgIJq/NIzq9JwrT
mmg2XL7eiP5xSRGhRO6dg5aDlf2lxyJRxnmQLkfy0dENuDKFaf2R8KEjHCeEFOP8n+rfMzJBkyOV
BJO21sb0JvwwN83Qfwlw59wIo7DuRSpSBEaZcMNMuOzhC6O0hH/1ayfcOll8pO6fAqjF01U1j0Xi
xZc3ZJPiZ5iDdG3i60sDdapXyxgX+MGgSxasYEc6usCaZBsXqi084WTDrxtg5vJjUCMl5ZvWU59u
RI+o8Goz0wf7Fy7klzjdSy0hruf9EF7Uplw+65ehvvmT8k2voesq2eFkaQgdI6qQaXUYV8bwSKoR
RXo1U8zarUVSkog5hP/kxzjG+9sktq2zz9ytP+NTQc/e3xM27N676KK+0wQo3yejllT6TTZRTRH4
QrPgL9jqHw0Ug7++DrQLmnibFmVyYmuiLleFjElgBwKgru33LN6YmG79gbZH1Hm63LEQbsRLiNWQ
GtrvFhDTp24VfS1Kw6eWepsv1z+0psnUNoPcI8HnzPK3uTZeRmrDgbvUZn460CCSZYC3qpn+bbhy
ixu/bkPsN7HDvcJow/TkWZ17kB3kFhBamvKmNCmgrM1y16ez1xTWUbYrCcddXhfFkBOHYT6saWfN
xRr4EdvTv8zct4JNt4D6yU6VDusw2Z4y2uEtHbbVmVZHEd3luEVSK0dePz2furirdD0cLvRCKITR
h+33/4nVqq7Fsw4t+2dde60Jl4nKZXbH0chewemfoHp9qc/ZQKiMHzJZ3m/v9kq1jmzBqqZrqETW
tF47R+RVPo/+Fn3zOaI01cyfAua4P+WWXkTVPc0EEqmXIq8bqHcRl5HFsLoCGTHbnQh5okcSfp/q
0YyquEj6WMYDUJlM1PtE3n3IytZWzujXAsI+NOerWcoYoeBcmQjU7hf6Hc8dLEykrzgU5CF8DWWe
mAv/ZBbod/pMEoH++e2tFqxVpCT4YJbrUIAfBOld2qV7/lLaM7AHLDnXTtt28qDEBFN3PZWYboER
aIyfqwiztyxfGU3UeYXibjgPAAI3FObT+Tlmd/qcRIZyudr+y7hME7hF+wXifkgGls3nPVLw/qjD
n30BVTwu4zh3BwL5r0EF+rpFIJoGjVzQlGyDxfnJh7yGl9QFk6dm706NXUDuku5O+fYE323JumbG
kJyowwjBoJcWV2RNeUOGdDteJjv+8tKwPlkU7HlAbdb9oVPVZb/rS9vOTbdrfAHl0kMejSXhNnam
6mCV34OrFtJzE0g/bP/5PoEjKtEK3wTrCzEWng/jwjFh8G3HWw3IpIddo7MPYGacSbMBzqKdn8Rk
vGC2TZLzIiYPs9pW14iPVyNJ60N2KWIVFJMT9eRx9Uj0ZVSLd+4UYaPuy5ZZH6wnQMnYmqsMbJNI
nja5R7oxToH143qB/gZj8QORDKyJG+r7HxMa1oB2nGJifEU9ychA33YilXiLKDoCQB7Fh88/99l7
LoNWsxdxlM9zi4CnltWiP4f5HAABHfULUqKXi69pRiiS7GE4jS6HYoNHf/8qpi78iFfoO70aQqIw
uJIiqk6SEBKPG6U+SpiDr9lI1Kx/FlXFRjfTHAkRANKK3mA6xs/eVGe1VEWt3y+j5KUz10I6uM6x
G/w33aHj6nYMuWJSIBxsuydfPX2K5zrfk0bYZC7IvO2dQ5LTHMJ2Ll+UK6e3Gshyx3+qDkZlu83z
wwgCVzBF7LZ1OnvVSNTYT2/d2FojTpXLELeHvigcA4QYB9P+GhnitDxfRGzkyyFh7m6dLTrJ0SzA
6A5Rn08m6D3gaSmdY+lRZ0YSsV1as3PWOj391QZySOgcjvnFP+vJyi0vygmDsaHWtMHJiCtjZ66K
ZEt+cUAgl9SIzHYLAtRAs3K39KgwJ46CNafCvEZhCBs+RfKQ6iATUc0+guaZWQAmMPfOjNGlaBFs
6dqjyOY56A2NHb9Azm08x9cJ4N9yhlGWY2dn5Lvw+va1lKo2neILZdekpIW5YIc2hoPzDXON9/SL
z0S/TAYbByBUubRC5HvCwkZ3UBWC0NQYsve9VDYXwMDOdc9FGxn3qKdnp/9gjHi/1Ctu/bTDKMJl
5I0LlYdd54cZkhktFQJoE4hjn41ctrq4xhAMhU7Sil+zltu/PwS4N0kMtmH1Q9q7TFTVT2YDqlq9
17z7caNAS+tKOyq0N85YJtYC0iTDFS8jHcu3a1i+DyEB0mSNSMjOUfJwf41fM4GZLpVbniI0iBeS
egE7O3XTpYd1lXOZ6u0OcY2e/VF/rErWI4zpTq2XZXURnpvVXxyGKym0AtbYuwkhw4LQUpA5/orp
EyCjVkRijkf5uxJhHFMOlTUlt/llh6w4c4AvbLAgfnI2m29v3QGbemw9npapK4LSwF5ZnchGEzxP
AKB4xPDoiVS5jB1lW5Cse8uWLcSd0K5176gIBsb8ASoEnmn1nLmWxgqfy0FeuHWL1boKOZA1KO8+
0bpHcVYIbAWq8fgZ8dEGpxxg/2e5tA/yEVYFhV3kllHP499ht0Dn53DhUxnVngj+6sQ90p0cvkgS
vFFwzeDBSn6lIZXL/goLnqvgLpI88e9Qao65Kz0B8FqO4Jc6I72ZEc1jEw+/RIsfAervM95Phlb1
6cD7BSk1wD/2AB818m7T+YNP/TqFzkGq3BGmdkKeOcFUrXHR4kGO8A+C0QfueP3zK+tpSDMMRvrY
sXS9oC9q1EOqOF2jLhEccaTPZLMtev7ANqFDSg8TkQQhRdjV+PflnB4vS9AM4fmlz7GZD6R8Bgh3
8NJXhX6A3Fn8Jnzcse2dNG0cXABk8MVFnlLsZF7DP+YGqDTnMp8bBvx+6AHtKAyaYvlOYL93NAGq
F/MyUZ3okWxTPVOfaUDAYurBBKq7iyRUMIB+RRa5MmY8r74U0bbVio7Qztg9FBTUA1UJDkOtO2iC
6JwT4tNXr3s2PozTimhuWogk8xgb4D4c/fo2bwza1OVOQO+v1ZSBoyp1vQYy9SQM1J8d1RUfFqoC
0FkPfc33TH9r7cJxk66yBJKKyE4bM1NwbQn5VqMUD6vq4sGomKLhAU6zTbPp8KsgE3GOys1jtrWV
OYLCc7x8r3/ZyyNPcKjUVCKrQTzQ0aqxTrm02fiYZCGFy/ltUkj+LGNkrpT+HTpt394uFKmbanKz
Sr/iisJ34oetjrFkODLgTwyeo6lnLzG/b/a74oYz9fYHWDzaxwal04UdzN/ozsBNhQgBbJ6aMUT3
3rn6JBAtFM9KpueD6+GqOUBGMYPmbnEDt6QtUtnj5HNxCJmMk7gpkDmOYu/Z0Qe5G1wwTSG1X8pC
Kqgawj0w6QgVCvYcOV+XUTk+BnNHJIfhhZVhpzAlYp5X2ha+SHeY8HZ+7Wt/ir0jXdXRnR4nKqFY
eKfNrQT5YpcPeoCRJkED8nxKpTCP3kVPl0qQEq4k9/Byw0qbgmZqbaJFOhYXSCZ/CYgXhl1dYNJh
VcvIWV8twnGaTGuNq2yYC32FxYD1WHbdxxCx0sIOsUhaRTW0KR5c0g7yyCkFOcYzQZkK9zqisyKq
06lrDeTDHf4Nqicczpv+fWYuxzqTeAkpSizHd/H6xriLvllcJEhOXMpvq5GSCp/p12B5feyIzgZ4
std+XEFuHhJFvei8pKJbCrxN026+BwLdwM1r2df2xOTIFBvHSUFn8/0lnZ9nUDEn7lglIdGHBY7L
1QKhItL0LW9SkLGJ64voFkpTQs0Jzfwz2win7WM/F9q7CR3hMjBKfW/DLUQgRaN7+cJQJLjeYD6e
+vbAGEso/LB/VQWY3W00cq9HBi+7vhWnPVhkeK7rUuKU6SW9PHaWvhDXoiSD9V19rbvDE8HXWv9i
URS9MEQ0Xcyc2PfJV2X4KvXvmc7ECMeew81xXRWzBoNUFUK8vjKA64rq7iyYuBEfBgIxMfc3kbrh
7LZGsre+KArBqtPH6Ni3+1iTTopwF/JcxnsXkG5x2ZBJ3Rr1g4Dk4T8ePv3PDWhdX9V07/vAsnCT
/KVURmhs7zc+HU8K8jIGydBK71XnxdFBHRLsU7LtvnbhIisblFmkjdyq86c5hkAmfucV4/NiFfVJ
+qptI9npzE3IzAX2PCJePGUo6ONSOhx/E3ose7nh0cGf3NOnYxTnaAcutQw3dfYSDor66cqChEw9
L0DzYrsd9Wgw1YgDYgaqvLmhcm/QJZ6K1LQuJAAkj5oW7dLfRYoBVh2HG7R67eQEPpF/8K53eQaZ
LlESAdoJ8Z5oZ3YndYC0rAEGW8BTWEZiD7piDgXa2gOzdY4AJCOJ1WsmbASk7RiJmk8bhY1h+bQh
IFcOuJDrBj+fBj4fBdRUckRVb8AOThA7Mc2ef8j34tx7SlP945aUMdZn/elDEKc219CbNG06DOBu
QfHlLQfv8UGMxvJuYpC5TjKICggn+Js/7Nc9UBG6NHMm0n1CcmrzUvjuAgjSGWAdyBJ5LHycsubg
MSsWc2+CDHIPeHtUEt9v7w0PRBGkCSLVw09VBI8pRpH+3peWbrM8H9cUdt5fDrSBlKBGCcedmtDu
lH3605IUkY/1VEthAI9VIiZ9omjyqKTx+D42RUXJkBYBC/0118FnHRn8mNVj8Er5zZ+9b7i0+x06
lgCMs6S/EdUU+SXV7uRTHDW84IH28D7w29++BcAJPweDzYscL4h3GuntnaD2rqw8E4e1T7c/6hyh
WxogzcwWZdwEehVFfwefmfiFe8vKY+oLUJCjHt5JcwX04B+NhqC89aHSm1MrwqonYcZ6J6tncP+P
ja10ckFeh3WimFyGz1vRZXYv5qyrvvmruz6jIPioyT5YANmEvCFDyYo1lJ4CtyAXQTSKGRJKHepw
3UMXINBXEGR1b4eX58JRNTTbk1vY3BcESwrJ5x6b6KnHcrJ4mf4FiRUzMd5TLmLPGJtJQqYv9FJ7
Fqj68iP6i0IU5X3DMsqBYIdBdr1C7kMZ7Rmtl4p0IQHKQfKFxdVMWKi3Zr3ubZArj/3WTzwi+5VM
nNasNnoxhbwN7vwiRkI+CwZbP/lH5Fzggq8sWVYEPNF7xTolToHRbSOzeNz58bsgm62yi1v11NVp
vQ3E+VUZixZzSTCFxL1cLmsNHqbxKn6gCNZHCEZ+JdGBAr8MOpAafgH+818Q1672fSDdgqzA/xUW
a7Il6IMAOfP0/xbLtStNawODr1lFOgMPI9m6Y8Ozuzp4bznFaOUXuoGp1F9NG63xa945KJMbtZVz
xLZal+RPTYEMo775h60lEu70fYqC4qwu7ANSzeJKnCGdNgHez+OL59Fo0oWNWIBRMhe1YiA2VfMA
KMtGxHLns0YV3AQ7I2W94k/gsVgoPcoY+eZO3BSb9CSMKoONIRHADj/WasVeiiTQr3yFxo6h5ZRv
lrpFA+ksYce9s8UxnVuA8SBnTWXcFE7++U0WvHWxERwFJhro7RNe1kjiXt9NxrG5HEB2yK/Kw7bz
tDcAJCrCUbMG2GaHgR5YNo06j8EzzC4iVBAOubYuxsE8JG/8JnaGaONrBg2dimdGPM/HaflsLHYC
6dKN2kmziAyJ1c+DCJu+QVRzu9caep9dlDgJwpznYraUqDZWYdpciGqqOKdAZs0Z4tQFeuohtZ2n
ihD2tzNwPiDVf3UkMI2ymhjkLuupVRILGPBzcShVSuACLg7K+T6mYElmF1gBbH1/alQHpUDtKSDb
9O+V9N7DLjniZu6R2Iducbp2irkgEoLskzLkoGvVHkPANlGxJOgUPBzb9AwFwT+i9YAxklcb/UJm
EtLjIqgsgMnDoFdpsSIoK0IAUGKA8EhoGft5QB8i3EQUvmkWBaFvm/GqNlN86m3shUfsXkpzopZb
y7IwKu1rBm49QXHfFGe3Y3Qo2UWC6bDCFqvxMVsoZ2m5UD0U3Hyo8OuVXlPrAyE511A53bWx2UzJ
XRqYgrY12KgUCLG0BcAAteFZVgno+sD6S8d4Wx93LheSDIlEUJhZAWGLIFBLqiyPYIiagWTCE3yV
kzZxB0ohdH5bF1fe2dplXEDulg9sZJcdfH8BlUal4zSp+VLRr5GWToHiWUDuaTYo7NHxTNGK+JO5
PamA+OojyDPBCgAUyw/ARS8SSGqkwx9hTrnXMY74Ui4fvowwQapUjHTCUcbkcGHVFmphNgOwKEnN
PNduNiyukjtf+BFkFXEmP29s37pyMFlmUDMiqxgOcRJoPZ8t9KNWrf7zICyes3zhk+vb2ycLyMhF
hiD1z8MkFWAu5QYajlRMDJK0AQOPgClgaIf57D7H2qHDy+cKvqFUpxfOoP3zs+fMXmNOUMZaaErE
pcPcRm5YrS+nsU3vj6frO+N2kfM7tlT2HF/0QNu9CVyUbf69RECwisYi5WA8AHpJtrURUJlsY+o5
t3XN407rI5LLGMbiLpBsBnwn5jyrPhmy2d7MwwYSElYEAjC70DwdQdOgIWH38MZCD8W5e52++Fv7
gHI8gHTi+ETncO1re/tFknzpZzrgdVVfABOGNq1fIkyvSl/8d/huhMo+BUrD5mvLdrsOjF85b3r6
g98Q+VNB0qEF4tTf7HxanZLi8Yk1svpt2ntJEco5JhqalV0trzdEuv70RF74bmnSOyYZFcTB05UD
TvT9SmJp/EcmwKCNpsX8PHk6FOvhrhE0sDjsygH0BsYOCt0k16hASrlkXRgLlljGclRS/DisC4E5
UfWcL9IGeMzHidNWYqpHSG+hC8MDz1ctXONXouFZjDMQwmHvrAsgVmIv6QU13/WfU5/UzAQrgw0i
og4Nj4MZpnJpOMZtBL0TmmoUrk5tDuAXicpNBIW4UkincK7/GLT+95tiaLunl5b3s5X12wqMaFJS
NwMjBG5ulTlmyzU8Y5ayeXFSzVaxwmWUNPKv1VIw/nZY/SX6DT6TwRvOoH++oUyjeg1XBO3r8YGu
ILrwiDVldlObBiOFHDAY/Znq+xho6SkqfzAXN91TA3euO6+ZOfDlotdcEuUwuHUcZtTtGZJaY6KK
kE1hXjjC3QyRkQfSss/IY0q5W81QZAB9ndznCk17n1uy08I5PFn8wPsskG2vem4dMx1L4luxsqIw
mVPghuSVPFKA2+Es0FGZZACh+VlaO9JkWqy/47OgBImfUgyC/g5aY8jUIdW23NVZ6W8ZRoKI/844
U0aVeus2mWoEZRov2zmpX5DMDzdVUj4Zee5FiVpvoue/mmBzaQwi2cILJ15Rib2eCL4MdPuCPalg
BTpJp7kExf92VQ+OLcIQmuUG0SVw65NEFoDlYMBWKrUM5zg54WU/2EDrmZvOr5FWaWiDv/BttqVF
l1+kkemMOP70UPX8YytOeM3KQx4I4Y7edF93V2ASlCs5y+PY4nhXKyIjVJ2zuLUKOC0lPAas2Q10
weV/WsULakV+APYHRvBn94PNYycOoQXKAaRQ4pWLINh+E91gQtkxWkKJIbIJ9kO4xtv2RAZCFM6z
Mk8sBcICAHU7gx5Oi3Od+8ZtNqu94FkBfFU3DvHFFk7NsodWvdq+K0ndqPjgO4a5X5038dEFmwO6
23ErkDpS9eb0HzrhjNdvxBOFaH1yQZcqWjQOswP8gXOsSNSy00u4CcdO5sYzH9ALqPE80UDIwJJp
1I5/99BdxKchOavdqBUYFnogGPnZgYgXs6AXlQh8eBeFPHkPEMKmOrnqKJXNsIGpw0mIMZeJLgJH
w1juXAKe6BVmFJ6BhK+HmnrytmaaQoFlB1AJ1S5fzIkv3FTGDlqKNPRZ82flMso/rojMQPIlt6to
DX+VZOzuGJxJcdR5k1SBMukaDRpMPuHHgNk9OXd4qZL/ELITXXxqJcZkVbFdUbtTc7CGVbwuEHCt
cRE376G2AZ72O5kZF9fKUD9sE2CK8gh+TJ2h8Ry6F7OSnfvflIxRpCR9VzeS5XDo/cSGJt8ljAcm
ledZ5vAT59d2XJONFzkUI8cdxl2RgGgq+Cc8RakBh3K+D5Y2PIfn80PC1reI2YpaLZMB7buLzWPl
JzE0OxTxutkmTngPF25K4QvAv8XseVGw7B6pnJStS5/a7A0frQ/ecvVsUDq4xLhidVoAcGQ86yyM
lw/zxq/Zr9ih4O28eR7ewHRbU5Mty/FLci7FDSmYsQc3Ahij5zZ4uJyahdoAL5EgGS8pQi4Gk0w5
+cdgjvkIG2n79btP+QcHoZXUKgrlqVxEQ2Fer1+zS3UhUDoHFCOPBkz2DP4pDVr7hsHqwcqRC4fm
71HKhf3KcgjfgnvPwVJYpSOp/HX+sD0rAtmrySFVGXLCvGMOuCScjRfPp5q53AhrQx6LsbLxMbjG
8kaTszea1olLIKB+4H1+9IXBqcglOoNFtYfwbYHIRzTqfvpaexZ4KJzrLH2mme0JFQOYOSSB/Tjg
o7a6kLRhzzWyfjYmKhZZmXLZLUWm6irnU10eF2F9X0cVVscANmt3RMhfhLS+5i0cl6pD1IZ72Gx0
jIDc+WiRbqKsj0uBl2vXUHCuXGgE61b9Iacp3ojIrPikNkInnaSi9K3xFk9OHpyiL50byfgLb/8b
wvmN+1cWKdGVAPrhBGsknJYquOSA2SksvFQ+9RCt7+raprZ0K7pONFCq+Y9gayRiEgMMaM/n86Qc
t9cEO4Zp8gv5tfb52kLKQFFPCqMxMHt/itt0YI2BY9k6Z0cy5/gJrkdkU+opxg1rYYcxbWYWAtoN
ZPRUUQG6e6Mwv9bh/sfuLX0q4qajPx+BcaST2Lu0RxXMYkN76ZDSsY04BPZsInpsVg6Z2ZRNu7iH
Y6j5ALlLDTAQCPDVVRtHqkCR4y1vwLchcmn3tpmeCI5dYqhlqyTdBw2bfGzdt+yQywdpBhK0uxuA
H2wfarTlM3F7V0YPdqi2hTpyTCHvrAsWRUFk1qhHkdhufghY9iodsEH9mPe+6AQIbQYG1OuwmFjH
jbjLP5zYaCYGFOvX7Vw9m/hPe5x4haHLWdYiBmFLzQphgB16KvAmQ89KT8V2fd8qYQ53jA184pnn
C3T+s2GDCXIAAWkfYCCKZL39O6vEiJ5W69jSavh4p+UZrsyvcFOoID396S/aEedheCHANR3JlAZu
132uJYXafdfJLFU6UAYEn6twAwocWX2v7JAUd+bhvshynK7ozqYKWwiZbHwGB0xHWcRIGbnVQzbb
tDytcZUK1ykzf1Hvv+9LlBEctv7gk/Iv9UuA08o66TAiIo0VaibkAUPF/QBxkBpKUQNLuOlrx7uy
F/b6bkRgsnPahZziNhAXsoXO/86uNwRV/BkHRheP//uithW1pks8Pem4Md61aJir+7wPfgYi6O7M
H2TqPQZmJxCCVHzQh0tfGwD4yU5TQ409S6MIHjaX75VOdsDKKUPbBJkPc5ShVYdO/sp6Kx46i/VL
aUFnGkzsSHoh9DC5F+gp+oRp21HUHYoRSwsJ3iFpgx1iRyMiX9JvMmBjYL7Rl1S521LutxpOujCV
RNdIkOAdF81dRKTFX6AazaKcnsLoNIKNc7sznwIml+/iMfOdIFf/x2VHDnr/9M+p/PUKlTwmGuDw
ZWh/4H4VpCVYHWxYKDIBjf4t27eOKnvvcjMHBm0GF7H+TUMXEfv4S0SF8lqQdm3TuiDUs28iAW6b
wBlvV5kgTu89Ue0xwy0YzRPrzT4XQEVn8Y41aVnLpUbSKWZsnoe2qG1p6CDje6/9n9CHTyESih7I
v5TMtdPwlZiyMCLIxQ7Mib5pylvMNOLegEpfO+CwVh0u+l6Jdh2SL1BnXvqN/DhVStlLEPPf44Kq
oUIqUPAYJhSTE9AvSvDKgLkvyjr/xkPQhuSkq8ae7ayKXvvPj0HueU5xrR+IGSqJhi3jBLYzGvHY
vgBEv6d5Oe0rtKALVuCgGzY/iOT5z/aSMlidC0xZN9peGpDbMapx4ypcV5Bl3UQbNVvvvPLPenD6
ANZNdkWbEBP7bFuQ4dW4vRwlBYimsIFl566HUMMGN7wmOAL596Av2FqnqwU11+YjLfvpYcwEfaVc
cJtDDhwkgvSNsVBFeOXl+pSJu4eIiz9DNTiICvzudvGHS49KHqh5ZSkR7pQi1QRq/l6uzOYw6q+q
mtfDKT3LTM11Oi1iiNqyD6DcqEO2FU7iCEu3d5q9Lc2b02jwbyLOfRHNswOiz0/CNes0WF+JbZwE
zrpeCoBlMGJQXLkzRJJ8ypH3vcMbiihRDtC0gNMwm8xllkudB65Skji+xEgLyir9rksypz8cTH5p
zCpth4ZSK9jpHChDwGijyScs1Kp7V/nNekqwGbe62A83+kjde+fQyfOLbLuScSLf3nS22e9miYtO
nV8e6j8UdrSTYY+Pdg/4azNWRofvURM41aoeQ0Ah/MNNywHARMIxBFrvMBqqVfb7Plpwh5b8snnc
3V8SO2ETYICjFJvn8bn58v9OLo+g6ZUvHmp9ucMhuuWfmMeFEf0SmthL9PIDjQt8Gvw1cok6l24d
+K/HHQZj5xIPx8MN6L3CsOFoSW8s14D/DFFevWaGr5uLqJ9WTbuoGXlwnHzZAXw2i5+DiAB/C4fR
DQvgXo2Snzn9F6jlF0dULgNtI7K5bOJRiPjWxXXw5FI1uWMxx3USC4peIvow+WiqVp29X1NQRaSl
iiJXEKCZaUc4+nqPM9XQCOxAf38f06P0x3KRID7XKPOifTc7NRO58K91Pu36BZIjseid2V+dqTTI
+feGYW/ZwsNRGyARNo/YakvOz5amy4sVdlAfELI1Cpjg9LtZFbRmzDgV/vvOm2crjvFOSQ1hI/Bc
IAsUVfqXwd+VQ2zGe9QG9ONak9nIU6kyyDz/KtrTvrSSbuPVWJ3nzRad2HETBj97DfrqKi1WSETi
BQx08F6hANBXnXuFW+MUxNUC0vkmDWbuzsC0fScnHrSEcHBcman74EI9VUa9POFPtktzJIdrclpN
1Fk5e8CfVzhebIIO++M6TR8fVUU4JYGmH5Z2pR8brwzK5Uj28mv79jKjzXLojgNZgexkRZlcvknJ
8mpx1FAJhKfQAJr5J7GS6zAQknpk4UU2XICF5tIKZMyA+XAkk1lxJ7ofYUqWiUXr7zFrvKijv6Po
hZxz1UaMmnC0VXPw0hJ8ApKK1KiSOC0SBMGKcEg7jDZHtdV8lvee3YmU622pqJnmRzf9lzZ2j1sa
IfnE74QiMLB/sqMZtuzDpX4VlsIRr2SJbVYfPkSPrWHXL/8ZvhjWjx1/hPNvlLrCQ5LQqq45h/w8
VzWjHiKrbFKNASLXKTNmVhAX32v36QmIDeruPQvwce5D6nn6q6wLV4ToM4kYH7C/fo8gPWZJ9/Kv
qk46hsilJeiM9g6QXGYbh61I7irzME3fki7qMUNSQifDjAZ7tHDAC7tEfhEyy6QbLaW7L5P8C2sS
kRrcwLy9ylqxvxpCwmfwln8HMi/cLgrFJe7qmSlbF0Ec5oM5LXFwbo/6fOxKirrghmZpOpnLsts1
3V3/NY9mR5yOiPDT3wEgxcsOR8NA53cwTxg3X6M/6UKVRd/qBgomxMzXiIMK62zDSi/lXfB2cPgs
pJWU830JzGbqMG/cXy9RhK0kgCLpet3r+1CUW2IDawYFC4IGhKBdqcvgXnA7DhsZS8j0/OnP9aDm
ZnGCHXgY4+5zGJHFBWkBE76DVicxkz4sTVbaa469sOlScPOJ3FxRNXe+pC4GM2eI28p7L0xKBajr
QY/id0dGUULfHdztwyQtC/1ATaRxDZ+LsfqfZmXF3uFzkJtjdQ7e4dDdVzdG085bc3bNz/GqpvVY
AytSL8GkuZEh7Is2BxYaQg/5QDlMf2ZZnEtQJnqzGz+jMLbystM4q85laXmTa1z28uY6FI5hjf2w
OhkExLl2tSLdBJbo/mR8tXygTNIg+a5V4tStXyEazQ2p1xCLj2+xoyD3OrQjT3HX1zFo7hVi9H0j
/NgYKavywLcHSowKMtJM2zhsYbM/AIdvcAypY6FxgZOxIW1gU5dvSdEgItNCc0tbP6p4PaujHzLF
jrIn5zgBTFwCxZ++/Oy7WrW/DTFJCa1GV3rynLxBfa1ov3Ge//d/sWvn2r54MTTuaL377Zr4431j
/9oQ8bsKK4X9oDE0htuwfdMu/PmSdddb1rv2F2K4ReqanW0Uo71Fn9HP3sIsDR0UxsxNDLiA806b
z2vuj9C/oH3obmQ4RTNg3D4skp2mv9VQvLBLb6nUQCmz6PhIdFmjFkzqj66LcNuCnE5732gcg4Co
tdqR8iCPWc1mRk23W9u6hzwNJ9/IbOwCuxdMwqIVKDT6/YueJFsQ44wlWHtbrNHtrVYxy9Tpa6e1
RaJY/PilfKUqcmyrMe3+zCh2VslRBObFrC0TQ6hGtGb1lOTAQhwStP1ypDZqTrNRyugERKHEinOb
1o9/VBtDDty1mR9bMlKIg64zcu3Y754KOKfmPp/h7EvZWH2VWqqLoIrToFFh2EB9k2L+2DJ+ijr2
m2jdIEV6//B0iI5mMXaUaoZ//Uf/g62JcsOnZZQ0T/P6cet4WiiilTI5zEqJqPgI/MsbYp+H+pbh
NorrARMrvleem8h4N5yB0AUii7dPDeXaWxF4WNKggAKl2IKl+1ARUmZW/P9MmImd+wQRD792GS4F
WWiHNSPa1SvJaVxEosfedE6SR4StfNx/A+InOoAkwrBfyi+tmn7X9sAGce6nZKtyudOxg8OmLoi7
uHGgXG0iZbLAZzQrUehm3x8v+EAfsG8+88yfPt56lad/VAj5PUaN+mVut4f5Z+16DfZOQk+0UJZu
iU+2Amba5Jkr/D2rRAQ8/0epcIRVs5s2pUn8CJgjlLexc2LWxcntvfdX0lQLLKR4S2bQi2APxjU3
nnEnLQFOqkiapOxgUB8UL7RkIi32+pIAKkFtG7NKEtqi/6XWvN3mP7V/lSGSQGa5qcZ/xFupElti
qpzTojJBV5MvD5RN4bQoe/1sG9lTnfnAVMLmkP1HuE9Fuy020A02a556gXwv668vQKpoUgd1aHcz
QI6iog7TksKfmQhdwmtT5mXbBvN0h3QxC0paBvunqqQe0sknn+adaRI3Xkt7ztQrZ0AL2U549pzI
losaUWzjJHQNgaPe/pGqJPHD84ztAnmIRUyUWMqayxeqldMHMcBgMnaMDTW0uUVawGG2u4CO36mN
4YJDVprPCtH05ENS6a2mqqZ53BgwINGxNeDrNmvDUX4lGKFl0D/xGfvQdzAgmFHCqiDk0iHmZPeQ
nDQQw/ObMl3/iglrr9Ruj9hfD3ghMZo2rGDvsq+vBODtinRAAURbs7HDjx6dA+1QhLwZoUuy1Z+b
JjzF6BvCNVTPoTUUcNbrGHbwSIXYAA1nx74l82tqqPDcUSxxD2s3V1X+2xS/i5dVC2ijD3offXQf
nBbJSWz9A7n11klscpdsJU8qyRKZ7wZjPXU5IpQavN0UjZHt3e2Z6rWVDTDcBy4NHCIMihqQ+Eyo
XmiibLTB/O7A4yez57Td0mlEkWF3iFlFuCq4rXZrOpoEuI8aegtsvPufwGlhshe1q55JObhSHYN2
v0oVHvqfd3jy/oE9i/4r9yCzl7BjqpnyJw9mYL8N9CNYVuAfDKPPnymByqZTtwmWHBE6LRIO8fK4
rMoGmLpZ6ywRTXBQSlJDqKmU+REAOk8ZAopYgATgXcgInID9C8y0S5frEfzHKevNq/owHELC1Hdv
GhV7ryIHCFfBi6/Cn0wfxMUiEfkRYQWwpECK88wVy+OChGDGsOEtbu5bp4HV5bft2Df4H5gZSY8z
Ud62X/8dNBGHe2vIdftT6quc2n5lMaFIVxwIzF5LZNvDJl2plZD4UUTQ2BBy27XT/loUGXgLjdap
VHKkNnWPhLiE9rrAv8BkeA86cIeevJ+COPk9LQsmYvBM4qUyOTprCcn1cKDFedxhkaQms9XEFzSF
CG2OdYgzRCLmol/glbL5UcYVxyxMO0BLSG0XIbnuu2vktA6tfnvF3ePXBkHyYUD3uctGDhlwsyG0
AKvf0n4uRzMrs43XmwSQy+owaypR4MioX3LPCZsG7ZUxvGGKgIp+8NUISWTMfrTciCyX8lQyOdn4
uPO7cmaQ/IEm0gg7DZi1zbMAAWM6zma5GRYe2xel3nRgovFyNPfk+DZi+abidm3WFlxNv1CHfdVz
QoHCGcEy7r+q4NzQP9QN9qIaTG7CZQQGWQx6P25vqtftFJ81kDjg43Bf+4F+EPzu77/rcfXKwGF5
4LvLKI3SI5nakxmrcsAq5sq4oYXv9jHm8USy++BovhLZhZMS/QchA2RH9TkUIV/U5Pq6iwUoa5cV
j6J3+Z34fbbq6IyuFHBwoqfcA2DII1z9DyUf+6pA9kUq46e89NPqSzffkt9+pM3gcakS47TV87Uq
+0IF2AEs12iy9ExI240jveROO+1Rc9WaGLUBrIaFcL1rh3TSiDAwnXvjaRIZ/TshEQ805eXDutnB
U+tSvR3lkbmMi4ieyQhdr3qX1ZwsAiJ6EmdBoGQNC1il1JsNF1806P4q6cd2/Ux/tyZJdY8MSv0q
B99MjDtLY5Nyds2tdu36tXefaDOeTtfy3rJAp/rwXJibqHeJVs3bf5wNujDgArNER1/Nr8yFLfQO
xu+bv3sL/kOK178dSBaqnt2vGYJMfGLfdjkVPQcx1c+GovEmOEfKbM7y9WQBcKuMxNpP/qcnGQX9
2Bb6mAKKeCJFtuLH/aG0Vm7sBDFsXx1TwtJSCPsoNY6TkGllC/rXRW5Rbk2gAUDCxlbGg4Z9ymn/
EZPBScMCnh51XvuJTdsre5ZYGsC2ol6GKVUBLWEq8kBwfk4RdI0kAj4nIub1R9lDiEwh/UIRp9Ax
qYazHbqjCX/Wvf3DKWldKhTfCWx6cFhT8FaD6k6K+kz20vNO+KZEghu06I/rWVOf240bLE+6GDVJ
Wm5bBJUAJ2t0bcuYNjf9nPtFWGfKXFcOaXTcQFDDrgQ26xG0F8muxC++GApo2RKYhG45tPAoYm5G
ZgZB7cxKacdgvONgGxos0IpPb6f10MU9V+lTvhL8zYQTmt43Odnj0fD7Dl4nOUk9vNRwAz6zuVAj
W/1jwf6q9FSqaC86DclZpXvGjNsMhac9xqUaaqOzsCzBUJUe9lcrLp6B3JCmkLw+r3GkXsNsTGEh
/oFe2rHsjwgHoXEU6JnxJ0oCM7bG3bqNekJiPwu7Pxv9/j5R03Pni5PhiSHSI5eltGyVZXZBh7/g
JRdbKs5YuzhawNCOdMyHZbUTo8CGrL/eEMB8p2xB4uaX/feQBwPgcZE5jPM679d7WhvbBbdBNerO
4rCnwlol3/h51ETk7cXlfcKTANhqEcvtQutgR0Qw1EvLN8U80qEr1/jT6rwlcc21MjpBZGSDJdIO
ugspe8+YzyrgPgQrSB/ysvhV7H1XgZ/N6/oiGSyN4wU+/mBLcY+TD4KVBpIVWawXhxl0c1unC4mG
gVyoV07tJ9yt4DMob1h1f/Rl14w9Ny/YdvjXhxs0stgctLj4r3FPQFFH/U//iKsykYbWHMRg51Lm
gl/w9xybMwkkaDyZlj2eFnCUc99HoDqRcqA5WYNMO4uHvR/8Uo+dXmfWz1EIbATKH6EvLE5N7XpF
qyUBug3nTMlltRwWr2ilErAFLDq30/5Ku9AFM8na2SfvlOYgpDg9BJ5G762Yspg1cU51whmKk15f
Ue6MWiULfc5wh36m0zVNKfYaaEAB01V+dFqjT2/seves7m4dLKxAJi/33WVHHm3NxAhIbP3n5u42
O5SSfD2J8Tj/04L99tHuh7HA27y+mrt/icQ1xLKhaDQHVsixMfxWu/TDFSjD0Btw79Zst1ERb+P/
1x7IP57nYMK5THqahYcJBBYom0zcbS4DCVILmYrKwHl7WgLb3nUl8VFoltGzZfk9C4E2Latqqfef
i8OwNsZTpkhtEcW1Ht2fevynXaWk+mKX6rqi/OEZvqznzR/CZ7GEBLu+j//AM3YM3oRNU5Mxchuv
q34ae97XA8vyLn2xoLEHqpmM4gYI5lfAhX4yIyIK1VMqgT+5tr2Y3048Vkq/d9c9DJeCCMIDOjz5
FfocisD6WV5ul/gYDcgKCHB93f4+a9sYdCmtV1PRtbrER3Uw0ASEHcYWNeYAtwvfJQLMGna8hu7/
bJhP6Nc0yZTFbWXXay3wSr6OH4gNdFHKcaBhwblrXXrDYUMbXl1eM24ZA30Dc7IaZFAswsMKzgPn
Nd3HjWeockTxE90KHnh0bk2d96SBAV9XJTQTxj7Rw+d9YmHfssxvbPvwH0g7PjuhEWWWzds0g3kp
p5s+GNqt6SqWfGnUpu/DpvfHuvRm6yLiUUqj4/v6mnuGAOhBMhUMKM/lGj4yMe3PEw6Ey+eJygO+
oExpI1hIeMw/lDcZD14PYvi+qMH4ZnCLD6YlgUbKJLvlhqOslblyjjoXvliQYyAspmAj9UeHRdGL
SeIY8RHL0ldvI2yRBF7GAXv+zFuDS9eBzCJaenIfzsUhTCQyzJ9zviRQ/N9k7bN4Z4oGgvVawlKz
uPmVkEUBmLIscG3ldkOOwSqDfHwaK4ES/P65vYn84M5KTKFvc6sSPiDV9d/EskAU9Ygu7kPdOI44
pIQL6I4qWlJQ9YqyTEy4nNTIhBueJtmTd7jILS8Tm3JMEDBsD0LLgrnvhhJVltz0GJWdpu12Tt2J
NK5RsYpE2gb+XHA+pID7lFcuuwjPkIIYfLq+4bZpyjCTdfB4JSeII5TVc5KlTyuZiEBmkpHmoWBj
1hd+sN1rLpe3EdnXtB429Skc6RvmeHxHp3qwERrazMTPH2Q9wYeKe9A6wPRzqJNuw2jgQBtg3oRQ
+me/1cvMQH0zuyAfjbQHaJFId9z9/YFJ8/inXuNpcMhgNay+WPPY1lPUe3cZ+uOp0T/bPpVWVt58
2pXecGrKwo+F4dC+MP7QJODCemGQTrHnDNIb1RThaJ9boYJhJe9j0rQCRITDWqES13CTRu4Zjmad
uYxrWpgv7OnCXu3056OJ9xZB7ZjocrtoVk6WFUxxSN1mTzMm18w45qaco0osSwe+t30KF4yRJBwp
WGJHLTJUMI4IIPdf84W8TvKOm3cMg/rB0d5nPsnr1c2OfQYw8NVSuAaMDL4kSE+Az1D8uraGVb9l
VCbOeWKEQ5XJ8GK1oScdpewT1Fh4Auo5xWq9V3PTShnaUNNf5sF1Nw3FDYEicE7F4WLx7UzvF/Ub
rVXZ6sxsgejhawWC5xa9rUwn9pR6en8CdvJzWIAJJl8kBhCojWe+sgPwLevSDhnWzt3CP2/ieeZq
8Ou8k74BBx1T13AunyEZQo9RyD5FP2rMeCkFKDRdqZiC+6dBw4l+ckx7ztGd97lQ0qCX2QoNaxvD
JS5THMbqHHulyWcirI87/n52eLbkfRWXugBVXXKT+UieKQVDs9V8p+KsXOkRzJPdS9kti9d8tki/
kn3Zy3imT5QRzcp61sZkDNoOn6OMZcViPwE2uhSXF08ZMtjZQZMDNGWe0+MeUbfVHIE4tz/2WmxX
QxaiqHKezuchOUCar95KRGrOSX20LSo0BlzEyocgZUdEMBII5Z19V1NSBaFPtww5hN5pBJQa6DyU
VGOv5b+ex8JzsijDzGLb5GD7a549HmiGmBOfdgkS965WJMpfE1xrGX0NC+tZDqzP7UASgYOMWy9u
AStxTVnhGIBY7i906eOA+K9JkLYD2btfvXsFREudCHs1G7okuKP/gcL11no72BoSBNvtRfrpY1bS
iXGQH7kLf5DJSPZjwIGz8c7jNPvL9o9zPoVBJS47/3ZwRCRk28PVb5MQJlb+7yzjrfnhOgWyj/q4
hj/8K+1+gRQPj0FFScmnoSoFuu+A+5xVikXxZZxeu170hTecCeAY3b4v4ZfOeTfZfpf/CN1m5N+b
Ka3xYJAMnID2ElqxEk56SivZO9sBazezR/lvH2oTS4610i59dYvadXr7Y5ySbRkzxsypqD0m7oZP
INN9GmBQilXk68p25upoeAT74T0KwSKz+QjCl/Qdi3VlSWKUVJWOOl2biLNGZjXusI99H/y08zK7
2RfFm+eyY7xss7cvpguFDJ5jHsbXOtYkAR2FDOXHdX1YtIIeltbXw1p7Uy/MxTUBVJrbBnTPzcgu
p49WIz5edleodoG82WJj72BOnmscBQ0XZoC4rL2a2xRZ+6G0ZY0qwDfMZr2dEmUWa8cVD9Z0mJV1
ID9lAzXT+SFUTtdWcNQB7/INZSz5qaUjxD7H03QL9+UhA1bEz1FaXd+ITrvTVDs1NOnAigs91nhX
ADkJdIsjiHQPPmMouc5aY97ds9BrifYnm0G9PDPZhjX+f7wTjHd1oDo688vldDQw3ZiKJwuKLBS0
vgVscBOA9eEZJIRfkY4duL16magstFlMx1QAjkBsfmV6LlYmXNDoCRLadfPQn5BQMn9R7n2RfNWU
yIox1QfaxZk1tEMo8F7dUpIXFa1KuSQxijtZUBxxKdME0fRIykO+5472pGNJ65maxfgiLfMLDVrW
YO3eBUWm9WRWlFyi+wYEvnEIvrhl9F2hJxOCnnQ/9N74YS41rvzqNzyTrebNqjajnC7iZzaGzbge
GK2z9/CpSC475SymbomL4n++fxMv2gWVIJ5q3/1NQMm8UkWvp0TO3z2l5/awilZ9kSZH3j7khNKQ
heZiRIhKC08gkk6wVcMYnNwavUek3pSkkMF6PDjX2O7iKkQsVn+cIo/xAStchort/9ssvC/Q57XN
pGVVj7xQXl3ApYpN14ajAyUgFsAcc+lmMjCD8qeCkED2v9KGFf1ZK5001ED+zxZ+ZbZhHavcDPON
gDGR+ZtFhKU+0hB3Mm6Ai4wHz0IBkA/0ob2HsSYKRIBIC02vSGpLC1d4YVASP94vPUgEsIn8OQyR
lIp3Rj8aaWLjuNi1Jo3NOr+Qv2AYUqTerrWm8+cGzexpu6gO37mQZgZlgULEDW+6XxLeCyUzioNi
rOIi0O6Wm44B9CtDKp7Ih02Qz3GgL+ffozATFMcd1a3Mmhw6VeRKlVkRlhf3f1wQZn3WvZADd4jq
OrZM7KoH9jwGryd2AYhiF8HfWW8CRzLj7Xjy1gxLeRfTpRLdNYg2xznnckYHP9Is13nifd++ZWiD
U/vzkSaXGnUUuxKK7fGJice42WmWOlWGnZRpn1np8lumEVQOwj5bLs1lk2TRImVjbGXhzVIRlI5y
3o+ukcQwdJeg2UOjjuXfIB3XQbRwCfNa8zQWomPjGcfwHEQh0SqtoyNAeBtSOa0GtED0iU4ktbVy
bGAUjjH6aAePr+xuKMHFBFN8u3qy16l6P94mLl2y7o1Ka8n8i7kWFHkOPjkw1cAp7u82KrmvBRxo
Top7ZLt9fNQxKh106jN9vAE8UACXQbXLUtLYAAAYeEL8t+sf917CmLYMEjvJcdKam93wNXj2k0ON
1b8fEouDfaHA2Mi1wRnnv2avJn0zDbAACqrh/f5MLzH+S2sD5zOppscHmDOG1kl5740RbTqfmHOp
80eu6A3FuLjTgk+okrB2XI4mak7QybMcLD0cark0uRH1VBMlmnuHiCkZLgFvRdC+oy/VZHjw8zpr
WRmVCBPqyJ32K9L05avOJ85dkpzyjb1T/jr/JVs7di6V9sG0zLJjLBVJEr00Gd1uCgdXaO0cYGqL
ndNdSlaD2T+w1bywQJZfQ95yEc9Tl/r0Kwto/2W8oPS8IuilBtmLS7rrDQ8ZnT8GJ6Zou8D07X52
2civ1j8FqsHzCazHJje4kiRzDRR1VmXZVvCixmaQjZ7k90Gn3K+2d0G+WJ4XiqBIaqN6mHZ8+PPa
rcoVPdJjpgUl+TUs2FwXggeeFooj8w7HOTzWIGJPfbZkK1Diirw80lLU+lsnNvsg/eimYQfQuf56
6JOEDa8aJI14js6M/tyxAA1gy0qSPG1OsY2ym8sWcPZS/2dWRjordsZdLXBwTMd5dC3K50cdjl78
TruNXZUZQEJUUL24etQyotTpcOYfArnl6opBNTSAjHfd4k7PSwx1EYXd1T4NbzJvYGJiH/YkdX9h
cdUZEylorSF5sdmFf/wRRYZKK5HSbZeJorpVzhvCZ57K/CYApeHOwbDNe+3h99GOXQ+kdnru42Af
Wv/KEszOWctKtBH3ElclkH7EdEcwmZtnL5in2tMWZmdVJ73GD8aX27G9Yz5DaMzrgqDpMvFOIiQv
lVluCIACvwNwISITfTvgHNC0Eotvl9sPRY5eHCDIkiUJgBajpNKeg9BuFMohul41vxg4bbhZo+G7
mqXPZnPnd3dYBBNdq2O5g1wOFQHO9AO0KMwHCQRYQxTTcufmMBPTBwZLusM0RtaDPFrb2BJY87k6
YJXXPAE9EM19ok1PdesgIzr6g5vbokz2/4EFWL/jrM8YHHsfPjAjN5QwSH2fE1jsleHJnoHo6WB2
Sh9Xc1XbLBHHgBvpu2048dDAkhun8iZvI/4ZmfQDYwjLvcheHBpXxruz8kZgsL3gj4LRva4+YVpV
uvYgPl7yvJcyo1VSPVICg5MWIiF0RTG+0WVSYaawOtwcocwHyH0RWvTuDM+MbCA+KRSd6oTlKssa
Vb7cdWLFZ87uZhbONyP7EmU0zuWeacSAc5NFh73YZltRTgB7tMUeWXW7+sohvi2h73jVbI4DNpwl
Hz8rbv6LnrxcVaKchFha+9fM93hcWaOlaAKPx8n0xNgPAHVPo2/A0UG+PABMFKpZhX4Nq78MegfT
i3PIN/ntoMYyPDPMWbtJnJb7UpMvrlGzzh4C2XgCGJ/AX5/V9YzFzSXkqke0GfeOrR5xjq5E/JGU
2CQgdrV+r/XM/D2/ZIksfGsLKkHQlh/gJAG/wUGbwSWjlxB3wGX8hZzB73RNkP0/SlyZMcprla75
TVVbfieO74BkMo4/B/xVQ3vMHTQvfNlfLFPmLfJf7v9eQfcRccm6lc0Tx9nt4/P/vnnMw3dRg6ah
70rV+EPAjaCD1RuphyYXuf7lhhuCZMphhVFMSr7VXo7qECFxmaSF/dwx1jj6bK0fTaOxeyTziJxN
TJ7AYSJbSjD/GK+JhA+fDKuGRV9t+d9MG7Rh3zWkCK+jG3lBVi5lK9ys8Ac2mNupqwWo0UuXerFt
iFibsRStn9dkthFumCBTGqm5BXyYwzYd7f4OHkUy7l9q/2c/lDZ+KnikHPUfnj5Ugl+S8rKz0zVG
q4J05ciMgG/X2MbO7fIc0kI9NmbusvNw0DWMHlvHKivGhQEgrJwn53y4B5ozuR/1gsOrDtNfDoNr
8yEWX6kPIWGLhZKKlaherrAvHFuup9HSwPEUukaGlV/WFTnZcu7KMPxEUinLrF+IpvZuVMHG1z2N
mNFZzukoqCRTiBntPvyRXUVQWmy+52U4WGBorsmqyJY/ybDUHqX/cuTD5VTnO5RMMy5EWnte5Jzm
tKSGpmujd72Q0YN+Lb2zwLcIql7vkbl8p24SYdJf8W/7Byr5CM4nozMwz9oaW4rfRg5cbnfEDgu6
qxwmgT/K+01MgQBl7/xWMsSKUik88/0LwYhOEcYSnkculMJdPf3zTqoxyWwwRwPTzX4JLwlpFxCD
+O23Poqs2VEiDeZqfIrg1BSY5KjmqrDU0cCfRnNuzHfCy32/IzU6vs4v7fMO2Nj+BjUKJUY+9ZIt
bNwcX3LbeRFIHPKHumCooCvm6H/FbWOJsGvmX+HAe+tWX7UXW5KFqKzBabPXbVuXbvh6D4L3ojP3
WvfGR6OGiOU+h9JJQmbTeaC6tKQL79tSNFVqjmthcGGzGc1qKQRuG2ia8GqbQFeWQ7K+ZY8njFgT
2JZj1mfSoQXiEImWyPsZaaKXIdPGv3yWUE+96NKeaMbnx/k7ImCIiJUAU+kUdcg/Xx6H7ujnoezO
sQxseJbzW49LR+EC2CUh9PnRr6ZL4GcZOyqXtxk6IS1UVVn9tWqPGRr7E/p3aWBtgh3YVvajudEu
j/v4B1LKaJyU6u2h4cvp1F7zW2wapLTFutWz1Lu2qdfdPjaFs/laFNTa7Xt/vYXJZJLenuIAV3eh
T5ntCAZjGKTTyD6gyMTH6q4LHOGUcoC9y/5hXxCwYXTJb9BAg9/CkicrsXApxfwIe3JsAPp9dztt
SMTiyqTJJNj+eLWxA9fy00EVwmdOK91yP0NqxLO1IipGnimv1hg40t2wQdPlu4IhOvMkd0oBQdc1
lEKNvhPZvmE1n5nEINwF8AA5mqr3o43YI+/wBu+BbWtSBAmsDESGoKYZYuuJmK52PX+O9IZlzohw
TyAHk5aXbo/F2WdjJfJo6Vqqr068gRYEVc8HCoKc7hsnI/pz1KgfqgQ0W6djL37phq08fZDaqDNt
ZUti7TAyY+Uq3ky/AlyVSVS9T9B0IfNPmDZQcJiLLYdWbVQzpwu0Itxd02zlQT/qmsqGRkycV6v3
jsOC7eZzuKiDTX4xTR2uSkc0/ygbnH+LIRyFgzp7OTbZZFrL1kdA/okR9WXWwgGW6TrGsNSwXGbM
IV3iMAuzKyd1sxV9pvuPnxxKX5PDNVvywVCMeaGY6jI/upx3V2poRm5CaMMZ7MceWMvr+swXrEw8
jai2k8hRrNlRUheFQCYQiWSjt5Rx5w9QfrFKQFGekfzNSFUtu/Y2tEHjScTpFFAZK6iEEs9N+U/D
xZn53kk7RQLjXH9zIm0cG3HhinCueZsGtCipkubIl5VUwRinsCFt37nk6ev9wDNrqlnWn9zEyclP
4NtRkhTG2U5iuxbbOiLs2z35lsGBifWPGxI8KGVPsKvNWOiWspa6ozU8kkihhS1SM/UPbavnw1kN
1Te7S0aQDS0mVi878jQi0b4cpyVZ/967tBn6kfL5h6V66yKE6gcxGfCd6u8ogJTrUZuqNk9GOF5O
aHiQP33cUUdiYivX6u6F6ZsbHXNf/bw+vOmyMxO6mvcsCH1uX3lnstMlSTELLOe9Ra4xY1iPd4DD
I8g00NAVTxgY/mQcKCxAk8ZnIDnE58N11hh/Jxcg2llm1KoVZUOgr3LxPo3VSwAXaVV14AoukgbM
feJ12a0q1AQT48iQLXRJ3rtddE6xRCTlfQGULx1nnOipuUJ/8IGw7pUMYGSuuyZPsWkVGXRfN0f/
+HCjcGcTmgHxUOKdK9WwYxZ+HThx95kUXljJLo4fzRZSr6djeGadLhaLj0lHDYhGLBNVPjhuZ3OV
vXzK3vQG9QHOvzulVYRpP/2GZhLj+5sPXldxVfdnpk6oPrjLbsU2c/a/8ozn7o2N80KXjuEJ/Lro
SUPuZWe4g+E+0rqsFkd3EwuFJ/A0FamOL8FQSEu7dKmC+FKEmZxfUkyCWd4q0fPz4+WE5W+cuAQb
8kR+kfYbcxEs8oX3MjSkODPvuMgGEB3WLSBUeJlOZEgNb/Vl1ZEAo+vDhnexK6kVwpzjLNL1sd4u
BnQohXqa4dP+wGvwFpgerOqEb27pp52jHGr2uCtwL3x+J54B3fFligE0CV7ht2ANBoUuMZODorIP
E7ztug3lvQWmt5JOrdqcsABOvDzj0ixLupsLHBCxyl8XMFqMtaxeKMZWuqPLxTMXKslFyXuqRGW6
0SayoZuKrDvpY8jM8t2OjY2jHMd/jXLo7OQiCIud/KgVo9D1ptOAfP5fqKdSkW+Ipv06tQTCPeEM
8fc/aMY4vYrHSaL3z5uR+w2s2Z2r1s0ZBgtKA9sNFUN2Plbv7zowL08AahqZQduh5rjucUfV+kpu
rghHfllTgv7QuVCdk/YERfCRpGQ2nqyNt347oG0D+1LxlOmmLjQpx0W/ymo+7K3eRMolUSKArXrK
B+n9bAtlkBTHegLB40fcyXb7nOj4D6OVW4+nQfuCUdJ/k40L3vsy9J4bvLp1pgbIy0EB7WgoGIE6
c/M71fl981k3svu+gY0I7s9ay29HgOfZ9pRjtmwoOwq70375A61kza30HsXhoquGPv7v+Lxg1JgX
FEc7zDpDfSg+NnEtJZ1ArbJZ8iYF4SBnPQ8qwdduQYPim1+zkfcCkUA3WbRRgDySZdVYfW5ryGXW
lRJuj0H8ZAB4r3728ly47f9hc0DgxVJ1Q9t4Yr7m7PHz6vPld/NVCe6XSN6Dt1D4rUHyiUxRDzj3
uBjUqBciuA+UkMCsZrQqGhGCmxpxzJwhnC1nzW9nE8VqTDPSemO1v9NJ/loguIXynVuBVBWwi6Jd
pIX9yLUk6FkTsbY2OOvr7n9zFV6aKK4yeBBWtmh5opvrlPyqkHJV0yp2Cx0g2y0okVa1nRb/En1l
PcbThsGbTLjEsD0BsxKZeB1y/CUkObyhoq2vIVVia0xJzi8AFs2qB7O6qoOxo72vZTiinNil0JVu
NuYpy7NROXnen73f4RvsvhESR2EVRUbea2KQ5FxvbYhXnrtIhjpsnfA/djsmUx+WQ75bPRYXlI7T
WNvB42QwR29DCcFp0WygKU7iWMNPkx8CxOMWp7740qBcgxFSLrS1PebISoo8zK9dSFidMkxvaXLd
JH4O5IHyAWmRuPs5ynRgqTH+wzVVFLMr4qnrqfGxt2jQz9cXB1/p9RKwXlD5RuDX2rnECc8uKTIJ
XpdXYNhjraiW9sTei0QSSbOLcSkCcr/RfdJ0vVfGejTMvur9R7PRi0QXM6P/Ki5ecKuAwvGzMLhI
A73ctjmWO7Hg8vnIwc8iuoZVt2JezOlliFJ+OzkBVKHBt833kA9r0LSsIj45FYMa9SUqUeKmgFu0
/jFF3rSZtct6BJ84Qw6rYZuU/efnzbh3A8BLqBZ7A2XAmpSMQigIxYWcplYmzHY+FZ5qiV0O8fmi
FHB5XwgTjOy+4DH4QIia6f3A5PHMZrLBphRHX1iS2k8xsUNZ7idXJFPSxubmhBkVWA2RIy47enjO
dq8MQ3DhJKSEhws6M2YS5C+DVbEVHqojfwAqAuQaaZou0eRbdbtFyTSmY0aOXeXSGaZKs9k+KNH7
1qCWwMmeMhHF5PjRr43nyFVsjlxxoQQpntILL6fj41OxX5jbboG6hniSGLj5RDiqoNfWP/W+dMfA
jdd3n3lbtiUSG9BZIUHgVHUSsjpz4IDFb3YKVUJAQeT9UxduGzaqFQdOt/I4boVU++4yPJIwgoYN
O5WIB5T36aphizAd1SaJcD7c5o3HQVTVFt5P+0271rb2a+DLaA0fH8IBFf043c7NKtXyN6wE4AW2
gZN8WJaN/2eAGJGFuKi+ML1AEhqzcIy7WRTp9LeYRpkCaVa/H2ynwcmJO69N7BiqdaI8erW/btTq
8j979hCoNEqVasN7FGnhfTN1BtBzReKH1lvXyZohwf1f0dbQKs1dOcbZtl1pOu0uitBSZojhS+dh
LXORc+z3tDCvz7KhjEYk97qudMzYNjgDZ7bGS2N17ZkH7nIoDJk1SYOhZNIzK+2ZnnC5+0iHx0ZC
QqsqI7pfLz227/j8dvsqyKTqwui7l+c06Wzvd5YpQA7h9PV6VH2j+GsdC40zTZalmXLcGjVB/VAX
k2mKjzd2A481N1/WTUpJ8oiEL9ewkBev4Fzb4+d4UwKndVSIo9LV2gQ55/9wpnWSxqNwz1YTiB9o
Y4TrDLqeIukPdB57ZF/2+vdLkOkbzS9nB50JBEXan8JEX1eq6uxEtrq1+gu4ZWmDjbCpr8hjx/KQ
5Vrv0PXLYU2JeoNK+ROMVPtOCUGzj08fc7LEsPd2Go4Rg3s5+BycMZCorkA2n7icy6e15kC99XiW
3H25Wr+UbyjXVFL6ARMoJ8IrFT6sWzWN2aHR4wvE0HNFqED9qdUU0UPVBZwhmfK4IoSWKxNruWKL
Gij2ofCf08DfBTaPk0zB77mirQ21jAOShW1k8chTCBA7gaBhOeMf9nabSHxpQpMJhEsDFprSOaIK
ZDN+IDMXAfnGWQE365hbOdMELvz68zusXXCxUj4wUGTESHNG+qnukRgkYwHV/6umyHAAiq1IyIWZ
ldgdYW155Nc8WP3H1k0UhMiYo7XhqqBpfB4Ro63JCAkGlCps+kSZnTKj4XzSKjzMrpechdnk8RHg
XHNUcarUVVhJjvlqsWfnvv15cvUXNglk9pOSOXxNEb65qyrgKoDbwJ6rj45UMVZzVeLGE7KNFPKN
9CHp3qYVXjDtVfQWxAxY7i1GB2uUmClXcNaUxdgW0OsR/nSQL6sXRLW9udKKa7hamDVos/15trC0
VcXy5XP72JyeRK4J5goAPKmAOrBgdMGRM8WUbsUiXhVZHw+s/CVCNAhIVsaUYXbWWRF5AiKc4xg/
qA/Paavmey+rIcwxwTIGga0LYwnNGSGYYwqRcziLe48mQr6chNPXCa+3gYvkX4BWMzHS0vUGX6Rg
INdSzMiv39/g9hpqfy7ZdsF/r/HA+xziVJRFhHgyXnJ/WBTYK3pZV9eynYDukR5JVuM67wDgJUv9
NZxlydHOYSBFHBYNhcFHzYyOQ/LGI2+kV1FfStnkIfaVBqsGJN1Naka3CJ6tgiP+Id7VS18duP1S
ljqIxU+HjYIe8Gje3cYX2tQFWowUchbVK0Nd0PLDvwsdxzRh35IqdXA+4AvlE7Nucg3C4bRUP2PB
BtPgGIPnwdj+s8MMraPW+HiE4Of0Kh3pswg34xWB/yf4cPCVEdr3nn9yeGKoAlCIdGXvBcqnWoV9
yXLID13Xo4O/5A9Wu3CycQPlqHp15zJA2onghMurz12cC0RO3Kqd9mrRcW6oO1rEdFdCjp8Op5m9
PVBWaTiizLNeuhkOlWY6gYrq5R1iQmZfHi+GS6uBF/oY3QcMN3QMOylPiQiRGYLGaNzGPwhaFiu8
yO0LPcxqx1GaIDpZT1dUHMwxVCBluEKM1FfEPcUaiXjUrZVBUDXkGp5ih3h9bLMJdqRmrAkDJvqd
VvcwReLQ5hiRr6xb1TDu2FPXM1BiqHMJu9nNamTx7s1j6stwKf2aU45s20uqIf2gJOGheU1xcP4Q
li9JGQl5DOEuNFRCc3psFb8BW7ocIHSFd0Az8gQcI4g7swtsP/XNoTWxZoRN/WSfyDDP7EbyjZ9O
o2153y3WSMekUy8wQOXcgqRdcya3qm1cQUS1/Qnl66urZJw+0g+7MF/YnKBpn3DZS4hgca4ENtwJ
oiaGk9VatvyVgBei/9jr83MhFKhA1cGn7YJKa9ujyhX19I9/lRVDijPvKko2qz6Osruh183DsTJ4
yARLwa1U+vS+5Y+AWsVkgQEkhbOA2I7wrJ6vwB2ieqZ84TRBarSKBaP+xV/kbj/zYWycHvDJ8x+U
jKZymph3dXs0MvBqs34ux7HrkulTxioqRFkVtzK8S1J5PvkgM8D9+3AprFfiVTkU86fEEJDU/Eb5
znLinpD8YgtWdY5FgHSIt6L3a82GjmS7z30MhRSgmYOGyWdE6fGCTnoYjaWXLFY8Cu1HhhCk3C0L
/2CW9mkzst9t0Ca3137P4Nnw8P3ojHW4dGT7I6Oo6WM22Slx1Tbp0odMiAfwozjE0/iFl2lrC2R1
WXTxtsJoCWWCpu1AD97HSG1mu/2Taf0BoDg6DZP4pmGgRJ7cqrT6AXV0hWvH9z8iL8oX4NnkVVHq
TXdXzsH+0j5gN9DorJi+ySoZiMb0ir7TGgAKTmiO5znShRkMxy3r8v3yRHCSshvRd20wp+s0hsbI
dldwH6n/JhUFoFf/DmzFbpnDuOP/9/EU3VQ/T/l+LFggycM5i52hWqBlaSEL4VLkCIyGBeJuIoq2
8Z7KrxBPVP8uYntfbt8vBMRTZ4hUah89ZnsVUrRhwCexn/rg+RczsmbP4l7E8PubK8kAouXbXZif
p/CbnPsH2IghCOh56wmdeaXQEpGald9mqG7I2R/GQKOsAUljTO8ojX/1JOW3rxxSzsE4joytRc/S
N2z2AdL95TfZOq9i6reVDY+aW/A3NkCADq0lmdI6dU3PUAk6V/5YE1QcM9Xd1Wg4BkTKpbCBaJiV
GdJAw7xstlzwg7GfBf1WDH05QVM4oYQnR4jOlOXY03CxQWfXd/cXQwsjYW1fGU76t/5QKXARRNme
YoIjKNp6fVoXbWVunOadaFdzFHte+RjXnKSEBOX/DRJHRTjaK5pLCY/uTq2T/JcXBWIn6HG6CKod
UzHaT0gD7euVIlQF07+D28ZaKnDn/QWzHlUm/n1B0JqwNylSuqqqSNR/KPZVT0RtP9z/nsLGm5Uz
Q12QyHrvOSlB7LVmn8CS6CCl+mlGXjrARlB6CnPzLdltwmlKaX4RAo9aCHcjGbS0PfvJKf2Oy1Qb
DZZdWmlabdUKMjYbmotktEzsKxLqszgDUTTCFP7yKS4Q764sxNvEdEg9p98ZfrvEiBYyEI+lAeYI
j8Pn5M5N81NZy0P2NCYgYd77G9EKeT1AkT3qvSqhdmS6unY1NjAqREn7GPjrDSOGbvCt5A3OGGO6
pCMwhIDuGmpms3WG/MJvMarclWitIF+vt9K7lbLmel4nAjjV8E6hfRXhbBrB5WShp18oxqbQzWhZ
U694C7I2s+VXEutvu3ov5dWLsjwMpJbGiVsFNZ6h++w+SmpiqwHLPUPothf8OYdumHYUEsWxrGb7
QKK0JQzs++puR7L6unP4oxUXSx34kmKgodJYdedLq7wHI9GuC9jkdOTveEb+1orqYvnhTaKP8md/
4sEbcw2IKpBPqD3SRvCrsM7Jh0uAaC2nMyt3ttSl3PjraYCbh2veo2NqHoqpl1LvVPyuHJZLUoLb
so67XOa/8LZq3CnCTQor2Z9dTss79xgqq7abo5ZvJRaF8RmXhgo5gOWh6kUop7IMBj0uFfaQ+rE1
uighEhEXfceOZsC3HTa8R/xODqqYHP1ruDszAItTXfQy6boefu5enBHgrAqxvExOhbUOOd0MiSaO
MZNsJA59Hnry4VEcAdS4mZYmeLb0+DKuCnyUFMiResRAcY9P/nQtuZ5HUxavIGqCGqFGzdC6Iw2h
sWry8tGVa/xpnUaMWIk4ealCbmyz6Y3HHOrM0RDg+suVJoPI26hvl1wrABfzGfB+/l9jXgZfnOh4
fipsiZ2gQa6jw8YGDXYOOhwpaa5IvjXapzZrwi5vhh14SDcQwpLLFenk+5dBe5RTGbZ/clbm1csX
KV3g4ONXHaOWTDaVl4b8Aoxxz3pBcGGt561KLh81WPT4/rwHdwFvEf01bQf1mM36sV8Cvv4MXkT2
js7cCA4zjldbL2kZndmFyozF0bOPWd3Y4g5Jd8vKoK5qmhnCw0lbevL/xQZApOr0hSAAkjTb2bBl
HvQ5gsmSZAtFbKkfkaT920skmxGJNIewqXpBIRvXkgC4d+1tlThWELZ4DA6HlUFUj76ArWIuDpPW
DzTjgMGdlKfIF5+7deEGxBSGXiteijKn6XL6nMcN+eFGxaLRfpm2yUoJp2M3WAXs5+hxabnypYii
HdqE2UbKFx5i9oqxTrfMT14UNTiy+UhfJ83D4kEw/5mmOtLOJNqTt0nwvoWfa2SezsCrP9NpBF3H
mWFj2ov+ET1eqzGd/vY44cF/V/ZqWM++GjayM33cWvrCi6p+sbcabQOH6XLsATfE4iZ1ncku1yoY
kpivbsdK3uW1gzzxr3e5GFsu+GUgJCgg/cPks9X6SVwy6RaOi6cacWuoDMGxG6UEnT7PGhYfU4jR
7t107vTt0xrU9gy5Z/5Mdx3q+DEPzfBR8o2pK+ijmyKfDuyf145z74htN4zr/cslMuDgP3qkBLTL
K80TezTYt+CIwfgRkxw6tp+bYe2suoPf0QTknd5LD0cTO2WmDesV0oJ2rTUVkSrx2V3K7x/khNyO
l25nGd5WUBKwQxVJBu58a7qLVOkoagjpNFWa5Rd1MOsAvHtWqv0dynoSnHrGd9Dzv/cTDs/yFQw8
pQNFx0Su/f3o12cvETRGRXVehNQK+ksHP/BtUhg4ii9W1RL/kZ5KVr4FZuqRnaeCFeDRbJO2qqRP
Hp2ot2FlqOZht8FoDUZW7ivoxocZyt3DPYEruJVJbJIVNqeLGYRZbikAfBX9gTYwtsKt5ZIbbGL9
CQJ+eDyT/uVHvJCTRp8NYiZ6pZmMcBxMSUbOPIojJGCpZhM2PcaQgb9+GpA8j1QovDDTVG1KC9+X
yNTbHfy6oiK/fUmPhtxqpJCmGS5b0+UzMjZywB+NGR6jKWpGZWQOXhwN0PgYV1AgqPb2GyLjTDkA
tBwcXvEu6clzIaxW4fD7DcGZoWuStSReHnFd+ISiceCCJEH0PFx4MZ5rkPnbnXrEXxNfyJWJh+J8
uvtu27jZkeZYT7UEVL7/xR0cOeeKEhoAebP0YzIYY/0LUZqnTm11u8LglCAfWXx1TgrKFwCZ0sMA
xq8mgZ+JNrYUdepKgWaQNjJ7NkTmOmCvUFNEfZcY/v+5esL8NDIPsSuXx3u7uAeQq53UtDmYvilL
pSyQ2ztzUNz+KxPyb8DSSjvkJ3OA17T08EY5ryrM97d/tkfJ46I9IQ37Ua3TGE6En1y8OE+QKWh1
dT8ROAlF519Zm6tew2csfmk1CDu1GYbBJCpdQ7yM+yrELQso0gSLtIizFYlZSjZzIwN/mr5PPCwe
olqP98P/sbpC2N/Waw9ewMtKl7EMqBIafO8596bj5ast2NKrPAyyv0sXHM61h5ElrOCBlU+Pvwbk
oJbq3BuqLgLfgVNQ/cfnFXL5OH7j55DVmH4//S8qaEtaStQ1HsJgCq6tn7lO+poqdTKjLui9zq5j
WB0/yPe4R/fWXyYLrzcRNdIllJr2oOn8EWt+B/CgTdmgM5VmgIemCkJKvYHorzrkDPJkERleTk0u
DxwKM//pgWJ+lpYBZTeY9bRfJ5KyKJUTXQO065vF5OrGZQ4zai0tzadxMzfeJ6z6WyHtsioe8oOf
JPDjaT57H71u+MdTW/BW5FXEJDT600h4B8VVzgv4L43LAvJnVSmb1khozBj+OzgSL+u5m0WZ1dzO
2lQN7h+zxCYRinmzCRT51Pvk6wDiRl6wJv6sZ+gu1kBfbHmVuy6Xni4K7wrGDzZL8glgFPTPqGih
4Y0cozB8nz6QfJRpcEqhUUyLBhAJCp5LAn2XUXsm8qJavjmcSdsMTFGq6p2b9htXwgNE0i/ZM25w
U86RNRzi7dlqCJ36mvqBYLyXnZdpdgHFmhQdglo52k5tifmm+3T0k7uLeglMzGcra0RVorPN0O3Q
VMdfDEdJJVq/mTD6p9g7BmhdDH6cq3TwqS96hS5EMJ1IdVKn2oYSIVH47Tf2hTZkBieb0+EEq3Jv
y5anuSYg9dW6gPaZVSlIqtsLIWzUp8x0llfugdMQ3C4ACHyppAO52JNgjNStB+bSBQJATJ2dvry/
yOlZN1Acxl/6UQwcnhEBoTR9mw3hTzu6Oy3YUz0pzwLdyerLCEa1kS7wMfaBAaCP2i0o6Cj5seGO
V6zwmZf4MGfiSH0tMpMkSc64T2tPrNmO2F1MURb6v6J0MdLjzVJfasWaAvj7gQ3OQD/9vOZ8g3V0
DOAjJbjF443v1+Q6uSkaxEsyShqHig0Fjmjfx/Q0bIkdW2eK6Kj56C+99mOasLRuxCKPh8+sAu4R
UWulUl2uhYf+HyuXe3lBApj0zAdA+kKGY/jD65ZRBhWAwQntwklRg9FuIzPGKYSlnlM7HP69/8B+
Q9OtWIM0OZ//xEglrH4oPmnyV49LRZV09xcRoYoyOrZ2r7xxfY40qOno7Rt9AwnGNv6i4tv2ZQkG
gLRttCSAiBb4RwBkY96XisY1YYxNIy1Z82EgA8+rRYctZCOxKGqX48GXV+acI73eWRdoinmTRJ6o
3qytmZO4g8cYoHR7uYECd68Alp+n2g9cKwCIQqxdi4Ke71avm4txCBQ2sXEZx1tFfxoZipsbL4DZ
4QITKofPHDQXiSLXOxY4IrSoy9yKFiNZiKL18otOivdgdzBVB0Z1KL48fY8eJp/cM4ZQSeFY7mKL
32XvsGsVtxVMjJ1dE1gPNSeLg+Hsl/B4DxAsADwrCVDa7UEzsOMusMASFVRzfdXbe7vQzWYrhNtk
CXIEd5EM1QrpfKIJG2lH9QovSQp0edva8JRJzBZWqlU1Z5wVHa/OMJXh6tADYv5hZw2iMupxhDxY
O/E2FjilDd5bKrcsIBxqBlmiF2PRUspcTj76Q7Be7bFQjI8sl0UySe9wVwrxzQXirFyQQ3OCel5O
J/VEtxryvYKJivrdlYjHqPoCzMUWur5x0cO86LDAM4q0P9rfgzjdZVzZGDnv8repqHEdjhVeHzAv
EZ/3W9oxRGiK9Tu1JNwkSOlWULxSfk0+iQlU+eHV8LYv684EjdgTkJsr2ID6vChgPdU49SG8lsOY
scLL3fwZba7DVrxbkM9Tj/YZ2LRUOzuqMolfXRIR+YkkgEzITYH0Yz3GRZcF87+OqCtQifZBxokc
mdq+XB4mzdUUs02hJ5kLX0aoZtuDAjwVMnou3T2kKEd6jZOKaPdYOsTLVwFR9TWsJQFkNv8/lSQO
VTHU7PCSAicrhcfPKc66GrfwmeMeUQxlyUJAzCbO3Y7LBNucUSBc+V5+Cey7Eo0drNJWLxMwnJyr
NiSve1+tga2ZEgEAPMw1MYbHek3VyZgNQwnEcAdb+OEApsQpA7oSFrfKvRgTPA+n+a1/eXYzpuwD
WrYBTSbEey+f/dn968BuXdWbtx+gTgVb4R7sqXXzH3Xf/eFRU/+/RIJQLiEqPifgDoXUbQlzb44a
/BwkSnJ5QxJyN3f5czmjuaHSuC1/sPU1M7T/RR2TBlrRAqUstl19lAZEw/nUnZQmPO+Sc+lex0oM
k6crJvWgK9JGrzG3Rgny+KUdw3Cyqcc1/WhxCqTuEXoSKJ9ni1Wu0soI33tuJOLFIp4Nmim3aqA6
1nN9nQ8/rjcmh0rfMK6zveUsNXTVrtdaQ3n1GJ3bEprg4TBO/+I5YlSYi5T/shkNviGX8lfsMsU4
Stw/wHKB5EvJ8yUmS9raXqJ91T0rdWAnq5piivC2SykQ5F8xzihsLo0tJkAKk5OZ0j4XtaCp2qp9
qxg3t54tMc7PM7e0Zb+V756e4S44b7ggHuEj+ub3bvyk4XDA+PkPSN+BFeHBI8WaH+/D+B2wWGAX
mXEam9NnqvmtJesZ6AG6UPZo8LktMv6WjgbI9IqqIAA6VDAuyKvqp857n4BheoyPwUjSlTI8tDwZ
TJSs9v59cCPovDBMkKALu6mTeFVo0B/SgHqLMJ9G5ZNCljT4o9SWYL6EjP/QOLWDzRswaoq112ki
v2JWU/sPgT0BMYl0djiPB5vPXw5YOF6BDzyBukn7NxY01obtZWnAdQOmza6WQve4/KTgBXHz1xuG
xgd8iNE89SyozuVG1B8blvqO4yVDV0UTB3QKt9mOp1X4qNr8ZiQbcTquCgG1nhgAaxKPOkO9egMd
yf2XJ5il5Kx0aAO8GZrNLDKUcRivnYMskJrktykPUCsX+KC/gQPAsuEkti+HuNwPvL0mlJbpPSjc
BrsKi9kwE1Ue3nSX/1Mkt/LR6TLT598U158gyuFWJQtF2BifRqUqjmGSHeEoZicfjP+ypb5nMw8x
f34N2f9xwhvttVNwJMQkEjhbMDkwjtE90MFx3D8h8fA0j5NB+oLr9pHFkEdfK0qLhbTaxOAAuXZc
6Ikhfknx0lls89HBXkeuGwaD8rjifXX0rb3Rx0eUr6XoBuoDIH+gvJ/jv2SsHSgnzR5ikWDhgd8k
k/YoXQhGwyGPRGYo4UVQRZ+Llmw/ywPw8ZUWHHMvfNm63OLiZV8F+t06leGfgOQony97tlT7tSud
8EL9dUTgUpksJ1WgHqCQ7JpUcORN2ISHn2XvNRShKjKzTbGotRFmcyotEMzj2FdxRQv43konOUUX
aGtPjafo9FgcOV0vOH8ZYPNkju/+/ojjZBiDAdmQe23fJLU5+kbPVrTdqsdkTzUsmKkzNO0dLZxu
aoR3zWS8Q4+yd0Go3kWOBMblTVbLoogO0epPts/gAoyhKYH01OTwFvuBV5z7SxfYiWT4dfOp46Aw
zUCCdYWeSojeioQ0zML1lLEzyo1VYVvEZ9PQ062cPAsA8V3kZDa/32bmFn9+ALH7T6ydKwk8otr6
p0yOWNvFjNsvumxydKpLpAPS9J5Z/tmpvl/T4DTKt/vkgSxP3k4KeIDlr8C/6pCKoxlHVHzYy4fx
oSUYlqHo46q74nMeSbn5nOxOhOM6PHwwbz/+MJD2LfODQpZ6bkKD7V7ryDk2rd1pz2inxPk7MPMn
Y1HzaaKhdsLBDLUVznZ+RWweChfk1V4GUtkMAJvmkLRTY6fv/pqK9kkWieTyDqB/Sn8iYT0kuo+I
MQmG0u4ymxsXL5LvCzWmYh9OdIMcSx9dmfyKjd4PNvjCS/LLEvKu8MkZ/FsFjMpgumgbrvQKZ/Fb
4JD/14VYC8/Y+wfWFe5IrFt85p0e80lxNsTnkC6oOEiwWWyZo688Cipivy8fIEyehfCdYBwPg2Iq
VuMVEcDjx48xq8m6uFeO7bkOoMsBN704oR0z6IHTbU3fjj1RerhFZ52j5V40ZYRSjOUqb8L7ff/a
gi0FzpRV4i5Zy0unwhfUU2B3SN1q/hJ6UU5CqfcokwKfp+qQEO2GZdCg2SNMRBzH5Gqv7Ut20Zst
AZiDVO2hr78mcTVXrZNyd0UeMeIFWK/3gVYsojbA0o3ayHsyJ0q2ainoynqH3kjciq8ihOM6Ce7f
R6UNuY23ui29yrnYK6jBTyPWHYrWMvvL5dhiaD52nkwcnpD/LBjf1/CPnyc0xAK0JHNs52/VW4my
0Vo/d02TZZnlczGmER1dUvK7eEjZn6sq6wvoDYE53lMjMFYKs9RD5p3EAzoWNmHQzO1OTbOoznCy
hLS4arYdOmhckb/B0/3Z++oOBh5G0WIAYk6Oomi0EIFsOVmLC+Jz6Muug3dFOKq+5xo60JoS2r6l
P0YPZnC+mT7PGBwk10gy89lnjFJ4C7oRGEOC07mCmLLFT62W9ttF+GfY3/PIFLIyvxVEbrKuEstT
t49MUKEzoSk69DEglXn1MDpXmJZfZCZHXb+kM5O2ydKE0WBFE+s9lNpAUdgyCSqgEGn9LtGCtTgH
5cl7atYOJNc4D/GXx2z8EOA+vphERADRgUg7DvtyeUCnJkI+VYs85TLTgNiyH5BUxFS2N8C158rC
zBWrrQouGeWrBO2woSR1MJiovooqL5tOFPzN+rNfeYehLbh6InkUxHTXnt9VyR+2iYWDdV1/2+ak
Vu6BJ7zGaMN2lpPHFeeeJPo5+uNxqbRgJulYUSNwaHzvbkkMZkPicRFoW5Wd0drBwhz9THBZepGS
58hPDdv5vcXr/crEuH98REsJJVmLnKsBIggSNxJ8NWTY5/eOfRb4ScwvSkE0dzS3+q8deOvjiuXH
aiTbB9lsetRuWCYIS0PTOoqNdSGE/+VvuZk7tpAlvMISmayLibVy68bxU9yrwdpuOcOR6pUtGtXh
xjAqltGfmvgkMoncRgeW7g7wmx2cZs85gbjJ2RouvzUL6M86tNAiVmv95PJqnk8lBJYgYv2S/1cZ
vfgRrymPweyQEkkaDLzrqSYvw8LbC53hf5ThfDc7j/s5spwpI8TmoJEWtxapslQa8qttS+PvuUrY
tozzZCs5T+XAlPr7gqXGpaBzvOkSaLMZ6mrNmrVDcx/Qcc04D8bdzG8v+fSshmNnORDUUdrAH7CQ
TC3wjupJOIr7eyXa9ZyrX/6Lt2S21XzN+DeS+rP/MRPYeR1z5OFoZP4/kV6KjyC6PYBnhkuqUzzB
Z5cXV5+kFONc19qSzw0meAK+TTo61Od1j7mS1UEPZ3FOE/obS5LElJtWbZuldwwLX4eob2/mc1en
T8K61DXWfdST6sCFq2LrXKKylRcADTUHKJsRSrTpdWYdR0zA+0CsCsxQBO+1Ij3AlMU8dXPo+exC
xavvXdYQDqTVBfaSIHSFAUWBSpQIRVhSy6/PplPe2ddV/CkAx2DQao0eJR5ky1hyrdXzxrXmx7jR
WiCSLT372H7pW4NLxN8muwm9/AJf3F13NkAiVyIHByzEOpOO3xkSA/7Rh5K//ECXBKGYxdwklc77
ZO5wzTLO4UtjYNyBFG/2b8xu+sewmQ34Xf8aFNc+Nq9XCKPQE8tfJsx/+s5xQlzu8nQv/VYT9Gna
N7I3C0WFnvYYwBrVbsOjv6r6y1vkw1JWfaII54ufF1S5TgDTzyfxVB0euSksQXDtYWOX+cH3KIrh
L2ducHzniv5uRnfFOPk46nJUXzvWJPLkDz8HcnkFZZ+dywnK/J1czWynyA7P5WQ8FCToFq9XT8yE
Xj9dCM6q8Q7lcF6U0q1jy6hTDbU/mM9PKMJf/Z0Hmf8quYLcir4iYasmkMxCl9u7s7sy8+Crusar
Xcd3tcdMg1VvlW3CO1dmB6fNi1xYF3QmBTMN8FvC2PvQ3/pCLFcYuX/G32eMnw8YNfn8Y1hQTdBv
ne3WOq69AjfS8x/dEZEwHHd4Cg8nTLyu5PQCgOqqN6voglOz5A3LLwIgGbJKvNHgwE7s/hyRXj7E
ZhFOVNBI0xWyajYCY89JgGvoHNS2VUMkdsM98nk9sG3V0Q3kaQ+jOB27tKxvAi4Swaw4BhW3zy4R
tW7TxBTV365cenhSYvcf9E2leVzUuxHi83UY5S3K+fS09xsM8kuA/UUUdI2lxqHN5dX5Ynn9PNT8
KXh21aJPQxbQ2nV/8AMOizAr1K2/RyLtVVJChnNaSMcZOteK4QMwvt/4gb1dX1MZfJZewUpomBkM
Won/5bDN9ZEXNHpGFS83zQ+SgzoKiw9FputJbVuMLdThPtj+OHwIP6fZtZodVhGq6OQmaP3AnapX
vrdrwLzbLvf99PxPQm4KPEisDnRTspdLr30hj+u2TLuB4A3LdH6r/+N/zk3jB27HveKYGTOqEPJk
wYnV69TBodtVM66f1JrPnlzkhs/tI7j1vD1IgmErCihl4i9Gsk/shM+YGvnG82DGqnjE0rvQBRvm
A9PduFVpDBjRlKtDDgK/Vz2ThL4kCuHPQJZN9lgN/NgrxzRTamkNqCZpmQlausjhYoNj8LudYoPv
g2MKDbsMlqZ0vxPSr2sBdWq+twkCfocYTLD5B3RVwzj1cI+eyEcjvANXFvGlZhONGHFhVDeLYm3I
j1kZ4Y0XBiue7O28Gu0d/zheBjP51OskDJOtigIlN7r3JRwpqQVlxgfYaAdc3MAoFU36KZ/0YuTq
pX8z8l1w47xN6o9+FL1dA8T9U/H6YB1VoyKmUuyYD+Qyo6869RH/rIE/UxIzdxQyvBzZEWimt3hu
IDgl473gUGUljxnyXj1q+ZGOFLuz2rrJchwT8flS8XrsWIkr99JaIbCOW9+a+Wt5ZrT1EIoDgNr6
xYV+gFRvVxyJoDveXIE5rUBC/mpG24ZX9J1YUfZICNI89D7umAwPpy5ulmoRhGpBSdT+mlRC2M3c
H8zvUU8hcQdUT1lcxKdy/eTOn/OkJL6wp7OCwYWYotIKlPLR3AxbjC7oZTMrdK/+w2tWH1vIPTtm
OpHNd+VhZu/6AXDgbe9H7RkEchzDP4pZ59fh4q/+0lleyH9lymBxKMXrku01z/aoOH8Lqkc4VL71
FDuUs6xV0RKknhalZSOI6kYjpnGTU+lb2/ix5enV7swUn7EfKzb3VemWrc2Cojy5pyA5N41tzvZK
zI53mKqLJvJszU8Wr9P0lSP5xIwDoRbHfA7O+5OPP4HxeYTJdL6yeQ6bDHtdhep8BzvN8EIk+dCa
I3BFACsR+uo1QGK59mQt0NIB6hJdAxIUhj9DQDfez+qq1ahX2LuU+EZq0mBzUvfzXtfYEOusPIEe
gx+dpchlZzDAVObqHXzcKfSuGR2GzCT/3Ee4qO6d8zKm2pVmAO8D5DslMzNXVtVZ4au+RY+tENAy
c/QMXNJp/kTotN+w0X0ChUAvGe89KJk3xf2irbKpdAoZ0NxwcIR36qQrS8z6t+v60t2ewmyLP98L
hxGE8L98DgZIptqs86/hDhFL6v2VR4ET8X1lpsqA/FRga1c5JZZ9zbWXhQSoGsvNiXYBtk+DQ4sL
lA2vzV77Ivw8KxSFcRP7/V5uWgpTheUxXPvLJwAmjExnx89rkwOJcq1drcjqJ+QaAarArc0exfSB
eFMJ+Dmp9j0HPP9WbIRMwDE6zwnfYLnV5/FDLd6k359Ks5upQlEr4hk3/e9ku96SyqSuXxwCBWZy
PcEWI3iPMUMpcFmvsMIM7Is/X9O9HojtK+G2qPlpHToqVtf3QTYD1kIKZj+qyM8TbbmcLXWKECyc
Cb+QXL/972iYQvEWw2wf5qeAL8E30bKUj70CR7uzZFTB0LGqSmV1WHOPDZKQklxSAcSylTb563vX
Xr/a2xOqIKL/UZfhqeUfNk8LmZ0KwOWctMLxq3js2QRvrA6JjHfEH8Qb8BcRIkhv7WBp2GU8usC/
pqsmA49g9YLXU2Fksv4TQ5qY+3HJ3UOGL238YekT/UlA7eW5QMItW9COCcKT3spUGKee0XhsStio
DfnoNs50XFfl5LCBVm8QLU7VifVTDaHnNfQ1aT3o7+qvFZsD7SkvJNrAllUjt15DJrGDv4WeSuId
mrg+Ma2iJeeZN6wEOzEYtmr2xVBRSIGaKqeuvAw8ciQMGEyEMI+VefT9WrYO6TMSYss2hGVWkX4u
jt5FSsJ9Lq2sorT40LGewiBGz4DUT8Y+Cdvdx/Rb1Tk5PLWu6Zl46inPdn1fGcXse5MzwW9GFaDo
/V0H3niitDuM12T6f2RRVuJN0dsPWOSU17+Vra95hv9Hmz0WuXr71Bz2pWhhHP5iu0EqSiRsU1te
ZJmNooJBQhu4A+FEyGay2FPtF4+Q9cx+JjV5ljYIqss29V96Q/O/PVAF1ZlBpLu2xOQXehZua+4m
INbL18tuc/GQmjUpOfC5UycTEsVcYgpPgB8hQY1TpGCNGFKgFdFkK9/rC5w2Q2xHu2OUkvEIYEwS
OK658Mlo0ECDVTHaJMd3KMjW/7tefR8QxV7p0sGYZVM+5Isy13/x4e7stVTBgM2/iQ/aOP8xfr4I
Obi13PONXD5p8a7CW+n5rk3mNmK1Cgx4sBMp9ojy7fwzCVbscVzsNXI7bApfrqN5PfOfVNVthDKD
wUszpJ0VpOS7kMJgEHRCOkxX5Z0JvCbTWz5GJOuMULULGk06cThm8U7ZmMXkhqYCVEYNeqEj3ydR
s7Ody2tH2FTM2TvZZhQJRIQUHnEBnUbhvuGj3oWaJHkr7bObHmGxgbIz/a50zigRogVz/VX8/LV2
05/Wc0xWo1WPQ8rb768U5nIWh+WxVUDgjbQP9DglYK7ORzIPJQP1PWb2GZNXmwN/t84hhp4L7Wwl
ZwCC6gemz5yvnX25zAru7GKSYhzCXjMdtsai5/PFlW4F3KIawrm6RUrT0uI53v7aKBgLfZjWJz8f
5rxX4ry+m4qyqKrU5pJtT8ByBGC58apsnBsLo3t9ilz6QZ72ESD7zRQDV8qjUWD/JUppvkPTf07d
enjcBZO6rM6bO9h8Ev95J9xg8rC8FZowbGEqkZOOGRaocJVsfkMF4bIVv8+GCQ66vxAfy4gUoOGM
IXivS9pC7izvTRMpoO1YeDDkw9d/QQPSMr95EwF3dOgDqiqytNHexUC1YCq/zpHS59Am4kb2GbHL
pGFzuITAMpd/1Zzopgw/Z3o4uBsIS9ar+O4149zZuA8PW0lFLx+S/kIy/SHgpGIbcxuWd0ylS504
INKWbPPYjAGzRBvBVoxG5Sh1I1/HAXaf15eIJxEzgaHvzRDzfmkpXEXZlxmo//V3JYIjBFfX+NTY
+uVi0zjahb7vFGSHCVhomqKwu1kE9hDi2I9CyOh08YnXFoO0z7seCdkgVcD04+wsD1BXmQj2SuLQ
EHIBnIETT2NM3AxKZqxlE/uV3n2f6I6bjXRijAjMFKd27T33XAONNJsmJE3nk7zCk0vRysV3mBB+
cBo777AX7YPSME8ym/buF6PJwkfD0JIbe+lm6oep2UCo9QqHvGtDUyrYlnU8ta1LqcBx8mxVS0DD
4CkTvo3cuO8Hv8t+4kBgsKtOz5Hebc5loTv4I8WlP3fR+Uf/rYEPfTV4pRN8oIuVpfKAEU1Nkxw7
2Ae23+GApJdwr1WWdYWc9uxsR/EwYZmGe0i6LXJPOOCVJjwdV1x6q1eqTmeB7qd4h2EZUfvYZw5L
/8xZbd8chgPrw8VTU0ZU85EguYu+qpAYX3C62eo8TQZIDqRHA/wYfftwCv+o0meZ2wWJVSBV7/eO
7lEFr0ZD3W3NGwpVGLIj0dwjV2O0gY5clNxmj2YgQtVPli52MTsjUx3/m/U8Z88Dg9rg370ZhJkY
4GgdSrFylO5byKPfmaC3Dh66ltkp5nUGQEjEZsBKnUwpGQlr11hV8t54V44UauS78DZR+y/PYdHK
mUPFIY7xIw/9uJveVleVWbYLtVbeDr/lPOK2qYA9OJaL0McDhCIfr7JS0izb3djvhRqqqcCHaYM6
xUmulJuWoSorQczrL1pt7rCxT8R4J03WcLWUrOWfTNw5aKBY5h0BprMMk3tWBcj5RcGHAyVSkrCI
IZqCgprsBSKMPM/itm4fzwO7ub5ezmAqFDG/BsNfnNqc3y5wTb30b9UXK7I3RxOZzf+pV2nJ5cSm
eBbX8g5BcIAU2/UpShaPjoXOkza/zYmX20IP/3tb7Wtiwb2lgrO405cpNsiOE64whHcf/yiUvP70
9XBzdtSZRKUgJMjuBO3pUReWjpF2T/tmWmxJSSb1l7wb57WldEM2yFPAlRSlsC7fAasEMQ06Vwz+
XJPBsnUISm6UNSNfxnTNpRKuDXwxeFwujltk4qk+kIhgRtDFIDdyORuMvj3KKwI7yQ/6ikx1vJwP
BKOBbeYQGqclQ7oRfn098RObjROkr3w2uxfIPIMlU2FzaFSVVm3wMPJgacjY9gumA6y0b0eoA1DV
P9bjkHl8BjAMzOrFvdzGf2y8SzbzzaacBkQ0YjcEMzJH1hk2l8eI22ew+D2zbjd3dUxGUNihtO5b
rndw/DX542yFH9UuSsnZVk4tEq1VvHpFCuVv0Px+hmT4vlmIiQA95SlFxSEUrtiksiw/pGg2k5c8
O75XRjhdCmsDXkljngS+o/wCqdWr/La97ibdxY+PKULsKZRWFtCRbKIoLFKJLuFG4Aa0ga+HW2hj
daIWtJZJR74GATMhHr8EULFY8V7Vw+2KPYfka0rq+T9lYJW1GWd0NmLdsIofusucRxhj0PVywvN6
L3Qx2voVWkQuN438Vpv3jSvfv6onECdRM7xz0Zh80uJ/Jh9UT871hhDjIxZZzW9HtglxUQeoFOHN
HK7cRQR90lE2WvWgsha8TWCJQl7cScshVkb5ZU82BXE4+Wd9z8KeaCEEBquKktL9jTElsVHDBS6e
caK3NjLbkWxP1TET6/p181Mf23EPgAKbEzqQqPysK4t+uDbE4q8JH7uQoUXm8iw1TjBKJcTCf3Rg
NrNDupF4dhhxpP+6TtmaH56bZ7YxkhGCGTQP0YmcRLz0o0/opjAoSEz5FhuFcTbOFTnNhtxAanQ9
pujc7HSUPpA61yHV+h7pXq15sFbvFDoXaxFQ2IAvrYGCmkq+EeBrlJRGXJJPKQEjZG1sHYb2cNLC
zM5djlObdDbuQwz+818HzAveF1ym9XhmSOQuX64x8tX7+esHZZjBx+AMLnolXfu30qbRjono7+6g
u0mS0MPQ90ajNj1ZaaRwQeqNJZbg5Ma70wE5pC72XEdarc7gjlq38AOxi2Hdhq6t19V/gLakMjD4
9vqkPkyDp1SXxNkxg6Giao8/NNsdyT68a1XxgDFQo8OZJu3AMsRGHzon+qvL5AvokwX9SC2izB8Y
iHJmtKvxEErYVsrsKKgjKNvjhaLJjKBbvCmCo2uDGaD13b8UvcWJIHadLghyMKjaUHbFA6PvgrVh
26Cpz1z4EAspfKep7uzOBBCd7pD8kP2F5eOlaq/SUkyoCN2lw2b2m/r8iS4jrazF8/ZC7Y6zpPv9
lelZOmZtbBAdetCi5cd7Mo1bta/6/3+vwMWVJCYjlLE8kWRetuOXbgv1ds13ek0+QReP0GBWZWXH
1VdS0FrO3rz83AHVUXcSR8ao0lqBvG7CnnZ8IvKuzkDKjFh6XOad57LnPr4JOgwN7ylaXUqn3v5e
dhXZ6SlTT3cNEQ5dED27tcARO0rtuvncXCqSQLvqH97gYRfVw4djfRKyBDNkWMSKjcyP1nHpOZKx
PxgHuCktwOBsShLol/MKioR7RbTlnSXT5s/x2BUnfr4144DKsS5LkCVIKxvNAk4PrtO6Ey65PZUg
fz2L1QIrJEG0XeYAAw3bFwFwDMSxHk+dZIc5ym5smNvsfZ6n2Fmw/FOMKfUB2t8Uu+8VnCAEgJu+
1DvvtGFSw8IPawgpGNQRu2ITy5P+QMS2Qt0v4XdeNicmCVc4Tnek2uXkdJkszlyNUFQYOY/8bENQ
UCjZ1o01ZbwQ/R9UgCSGB3mAmnm74pCSJiSUYei/00NSA/W6HL8wLQM8XWtOj7eQCj6rp9B0jLQM
OftC4aTyGwrVXpnLpZO8nAj3UZZXtuxdx3jNShakAY7nTWueKXNee6CUyztW4mgsDARxvoEATYNo
4YqAGzFhIa0+hMJ4srh2lSxCJ4RB2bXfuU27Rqvk1om9l2l3LWop2EVKAyX3PdHtPqqPAxlJ3OMT
NCCAFk7PC5Hrrh8+/+yMkmwf/4qYdb7m2bIE3k4p5nOjYAp3mTqZXLw6ATbMfxEjf31DlWEk9oaS
GVqNcO0WLz5h+orY15Wrvomgo9evCDh4u2vu2lY27Hi1VV/RWlk9bckMxbNGFT0UQUDsHEkoGKDJ
nJ6xZGXtQq2FhKE9T67sNOR/++zEZ47XtQ/BG8usODosglbBX4CYPtjzt31tNDJAPNeyZifShYRC
SstBq0xvWUn9+82mupLfQUeX1GaXUBXNwW8YRHjWZkaxQdDtmQVW6aajwO2cwhzMHPIJXwwbxiV0
FxNn71mfxr0dcuK4Lc1UtsB4NB7pEteobuXVhHY/7pRSRYjco2AaMgwMT27rTzTJkLNT83xDs4Tf
IHz1jp0beYoVUsZMKaX5/eYlTCoxtX6Y9FJ5Vx6DOmYIlnj8RhJOakDIxXPDEsRuPTOa6JrpGszg
e6nHmWuSc6heQcAE0SQVQSePSw+XnVSwujhmzyuAaEWenqUaQS4z9I+LCmS/PskTnK9Jw6pA0gLz
BS5DfYL1tAJSZI5nyEK6fxMmCzXikN37WjetFamta6eU56dHTTLtE2VGtrwXgnbDCY8nLJBXZKRB
Xv0yT2ErkNZD2YfeuMxdjTwQmdBQw+ZgxnoM4goAXaKLqYEuNV9JWTQqlwIAPxWUK3AcOIl7xNUr
UCsI3MpI4ACIBEgOkhMzO0MGKTBpDDldpfDwc6WsEwjOee267ccjZ11CKAW4yjJFxh2atvGEzJci
WWVT1xaZgGodUjo3l+legrF618K7jkzSfKPszjmjfRS0NedzTUXlyjo4Ot4VWKPEU0i5LlxAtvqy
6EVXr28wAXUWzC7eWl1BpZeyWDUedT8dvtIYU8aSze8fV3z17Zm/sLmq7X+Sf0tglWnmBwT3dLup
LtW//y6n/sS61iJBsz+q4UraWXmifTaqjoeXdOJBS88kz7Dbktl9nQOugbDukSO0XRLpWLOTSE/l
ZdNCDUY1asRLelwBiQBOFWYp+aEfzLBjRoZnxHKWe7Wt1syMnq2en4BgDYSSb5VVRI3ImJzBycrX
SD/nwz+v3T21YhXM0WLCYXqDoznpCa/m8Qyst+ArhzW3+DUW6DtCSp58ttvMO6pDGnndKJfhGguT
EZOSvzr72/AI2KKW1fa3BvDY+pkCDRspTTzwDMpPLarm2LmHV0sjH2XXck2FKTO6nQ7C/MhQ1IqL
XJa0i4P8J7qCska6DMsFdVy3aCGJ5c3GPwSpcbzgZQ0KmP9RmB+FQHXxVmS6rYQrt1qYHYZASeex
k9gCgaRU2BS9PxCe3i3YuY//ccsWVLdHDh9yOeV6qVDi3HeKLCdWQEMrDf2PeqsN8YSOqLU2O6jF
edp3scJGRCKRPYEE9qlvpL+UDK5qSUnIs+MiKpMe0Z/HwEUCbDtlVtg/9j69bMfev9dsZvsXs8eK
gPBevJDQDJYWdmGvQeifpQUH9dAxz1eM8JR0JYabs2kl1HVJTHKicYQgOsgjmnTmcOY03HP1Ep/a
JNHtMPwTH4MGwIIhWRNLbhWx1LJt68MM6QKQ545VjLutLw23W9AR5EaWss2G7pS7Fk1d5RdPNV7s
xFBBMAEUXUSM3Gccbn4bmY1CMp0msDeM7YlLWpuvhxQ2Ks8ia/Qg8hO4mQOMW3rqmZ22KG8zb24o
68yShiSd+pXphp5BKAw0ary3y2g/+EiTguv9EwTBtVdk1nIwrwPDj4+HHEHB2r1BWNT5vIsngyL4
YXo7AzRZWJQjgaySvso4rjFJAQ5kdwd6LCfIZfwdJr+70T0N3cmSUiZzqeSimWi5p3zpELOhp15Q
OUeY+0G72D5YIWM2UJxKZn+mzxxU4Vfnot46F+g9IfjZYI0h44vc9hsIVA7yNZ72c7u8rUQtF7on
Gyiru5V8P6KV2q9KcvxRY4TVsom8GCDC4PIpQxTIvJWe9QTVKcC7sPNHz9SfKTQ+yo3h6xkPqNrG
wG+lXWyoOEDDUH/dbMgyVtwRNSr9hftE65wHHlYG9sAOhVI0QAmZvZDIJhvxCXGQQwqCI3IfGI9y
tmV18nY4yjYLRNsGEeeJlEc4CQaflPiOgwG/xRgPCAwDMsaQRhWNo7fmrqhBaGHloBtY7DHI74OE
3lzQZ948NJa/WhA009DSwLic9kKKU06qwrWpm3PApQlD/c6ddjVe9lBHsrn+n/cip5ijD5C5W709
gV1bEcyce5OzfOwqWOccWqjExYk43/LO/P6PTmm3A4PuMhYoBA1/cgdH1pqP1BoktwYxhWpk075Z
T1c3DoMitd9Ih8ibiBcOLw18PNJAGyGEUjuRnzQHSWaSQCYCjnJQImbIZwVka1xa9QDu6C760BWG
koOhykhCR/nD2jAgOTWKhzp1TU1Ou4VUrw7k729G6R+R6l9EyXn599Q11ZqT2Eta/drM/beHmO2v
3IR4VJBwPE0vFJWAFGOt6Dlnox96+AS+ur/6fBf/k2B1UJynWisBJvXu9dNyRMN0hvZNSHSPiGql
PbyL13aiJtCJIwad8A7EQd8/2l8t88gudQsTVbD88VOLQJDsKYSkFWFa0nelCc/LJnSWHok1w0fH
4GXzok0gBxvcH0p/G4luIF6m++cyVPmExdwJ35uXpMe2LpMFCRHoBEhue+B75qPo0E4CCCwG5SMW
jMQNf27xuB3+iy/eMx3xugifHUl9HrDVc/K9YyS7YKfk/mSin3ZsIz9TMa4Io1q0xstGqC2sAaA2
KEWdSHkzS7hIm833rhnjdvyr1JJ3m6gE7jlwBgVylpyLalAaVkjqhb5kty3NEhmXvVmnQnj9oTnt
WIthKlKYkZHqcHUqsdgl8dB5yA+ZQIurb1qsWbsC/N1KQVV4CbenXybOXaUBzu2frCzKx/4EL70N
fHIvI1TgJlw+S0ktjECyzK6QH+k9D92xBwyT70vJG0V0jbeo4s1nv6Bmxabi4+Sge8ewUKcDyjE+
bhdi244sU/dAT3WWEV5bAIm+KIKz/QhWfICTZj70Zs40KPT9NkWKHC2SdaUMsBmlObAnvH2zSzJj
nJj5+zmAamk8bm8XJu7J95tEt+B2ZmTG9JyRMAmvKNJzecHg0vkGphEvRuaHqW3PI7tVrMeoVCsq
QLbfz5jHr2msMyUPMYrO5yP2Z4mC46mZIQf8lIUrK8eHmKn2jlH/HiN2SaGnSq+afdmfuGw7FcMt
/FozcLvLmVOdMROsmuEo/0wgyIqeG8rQyGxo7yio+sP4dt9b1MT028VJiEc15qe1HTDS5c1wIXEy
tJybqaHJOsLqbwvvaxJBzgVXSwQrNwkwmrowXV6wREVhqWt3/F2M+ZFc6anEgsg+NCBQ7b3iKCtG
gKgAEAHYRNajDFxZR+kCxp7tzNa7AMvu/P3pIjPNOnZA+k2whlB2ILQxBUxbhwPlRMZ8cp0mT9rQ
Z6Wxj10qbuo3OuXRc9F9HZ2T/LGBie6+aZQ49MS3IBqxt32wZEEqMVKeoKpDEtKRB7ttFBi/j3I+
VIZrj6iLJR2uaYMkOKyIjudD6+FI4pIn83OBK897Hf48566dHmyE5D5cOme21YklfGYehOmgZeeJ
lyKp4r3hbhckAZBklGE9aS8iL3+Y9bsv3FH4zouUqvdpbBgrp/t1HSDoC6qhjqDoA5h5+02383Iv
IXSxaXhUWBUHQmiIkYTYol4J1k4Pfit0ukibrQAw/uKS/iTAbVwzBMFzKJjFLDITPlPFOxhTmLMX
36yREPzdNeElB7gNwMwwHI/BT8X2sy/GegROvo87tl6X0+wuhXpI35Oq3JGrZT26cYLEUlAxvC8z
AWUUC1NNua25WUBF4JxLetig8Uj2tLwL/HCoaybBBoXnMtQBbqRFMq3YyNW93XYdCu+GBAfWS6Lz
nIOJcBOOvbdR/Q6X363+KgUdnmhxSyQg7iby1/8fEuFOL32zjKml2UDTf9viCnmZ/UqRc2ulDb/E
PIGlZxUofW53n2u80GZWrdgUSv6/VGtPkl3sps2GqdtQ+5nSPFkSR7+dlm8uL8cGgMZx9zBdjf5z
a5i++NmlHkUmOFeJ9UCtwjYKrzyNB8ASqv0151MQ4LfYrbcsSuvNsjo8DN+LbDdiKUwHl2wLkQeT
ca5GiYRWUNbUidjn2/hGpRPFX4hp0vVoCZbakjOmLCdOon9hPBQDthYrgOySgEVrX9+hjnirdw/f
tUuO1EbwP0JS1Gye5jviSAW1qrPMC9+oj5p5OuS78c4j+SLrYWCg0pWohEhIdc5gTKJbYC5oJ5ir
4qCyK6yoFm8K0bpQwihO6rn93hm5LAwrTVJgXvNObR4cJMdFnGoZsenC9IdrwIQVD2yrG4co/VKs
lppGt7Ma2/G+dXoD4EUHnrdyGnb6FOJ5ImuEv2gFNOU192jljvPLP08xABnXFWdqKHzmYfeWv7wd
zL1lhfJTaNrg45oRSrqSlhkXqMRlAXWe2c3+YldR2qXMzc0b/kZ1g5BxIpwWWAuW2qAi5650V1Ss
WEhUlwibYbpxGapWvkOAfoDHwNNB8OqVZNshc8eaY8DemkfUbO0W8DvXk9JECgIShFC4iB8q5EjO
CuLGn1NLTtVK+96HvgP0SiSIvw0jV9FGGKNP2qPvN3O/xT2LZZol/+pEdfx40gw6RB4e4XBJUMGN
LbWYG9PL5z4EQLosvtocIdLf1MnH6LWgO6VIsnC+R+T8uKaJinaHjRc01N7/+WItEU+gTwiOPczP
ngc29cOoXaiX9QOu1fNxQ69uoN0SOxyMWdAG4X0ggOTcBOAH7EUoHOgmw7FrHgsBSHzjYpH/bxXP
X8iZCKXQUkod/ewI97mnnD19TilepOqftQqohlelnrO1OnXAAz6JdkZxRkI0XqCtCx4i3ORWocsO
GN3lV59lSKHyccn7bWPusBQx+xf9WitVGvuqWnf65MOdhJ9qCtyVvM3Fo/rgLQtqjyUfJr+AXGt6
5kl1JosAjumnnNRLeeaLlR2IBCkLuv1jSFeqPVtUxDnbT6yONHrjBn8cqbsV0MzsxQ+glyHdPvOM
ssJchAAeot7jBLtqLNGRgwElkGAxcBg3Tdl1fOujZ0HVf2IcQ+kWDbtHQ2WUZI8zWeH6NBDYrRP7
XqD+L1wazYWTxACn9h9DknTZ8xla5MaowPewvgzAazDSpcy40/4UF/ikXHH2daMV5divNEVuGFU2
ryZbX/QwbH4sD4Hn6DHjDtuUt4JOezgGtIhSmQ27eFhbNCA7uyubmttZ2gGuVS6fzkWTQVKaCpWc
Fu+y0zCJHJMOtwMXWkrzW8wiqg2FZTaOgU6RheqR/nfrwrCeIKjW9+HaswJG/NnpLRXXAjtz9SLd
xM9/MikPsdUPK6p46vX+G07sRKvaWcX3q4u0tSe8lx4by/P4zAPJRoUr023A1zonTfNTToZL7bbF
ukZyTkyNwiE7hbCbHnJLky0Ihd6dP5PRsSp7WF/87lR9nd2vicl/cV/yH81rYsOkZURvxqPuUuQZ
cC8I4M4MBdbS9yYj0yJ6W9m0Pn6A3/gkbRr+QjtB3XIN4ao8k2mgfLJOoJI7kWgQkkbbZ38e8BNe
3yY+uKh0HEjlhonCym9bd+sE8z9nSYSEiEggRCc+vEfWL208dV4ZkC1vwlnoe4qmlKgY/JcDZwsW
YCWVSewwAI1W6b855WWXUXH2GlMPb5NqC1ZvH1kWEJp0+Q3wyO8uxB6C1d0qUG4uJoBSNMKFoike
GCtRu7a7Lc1nAQ/gphGwv0ZTy7Z3Emo5K4GKAxWc70iVDYyWboLgMU1OcDmNO2y0Nypr+jFciv7d
2EZ4EzaA/hwCpcRKtAmtuXRFqtKJoZByHouV69fXTQEHJKTGiYR4LDIaaB7Ly/q3bdTWI2OC6RD8
AOtFUl6RpbDyjbDxFGcLtFhPg6DQQe/ESEFahOknhSP43SLrpahORywbksGDjt4Wot7YejuXFxw9
rkdRX+WcP3uGeM8++9bfTJHBxcvXcTpBImhAJjH0258PiVhge/6PAIP9578RC/jshQaMuUinc1bh
ryA8qeyAbK5S4GU97m1rfyKrZqvCbHzKjIcOSSDW1yH+fGcpRMhOODf7AJ5DlgzQUswCXdz/X8EL
ywQFiYKCmuzuWmlTN1+RseBoNOJiyhoQGVMuIz8AHNj52r9pNModAKuLOgItmfsmil9eX6LR9xkA
TdHhTAZwawa/b3veCc3Y/9yiJNUDixk4vZSyhSomU+gyFYCfiu24rgT9ym5PcZH+mWPGx+UcFL0C
i2TYxYAE0DEHkpIK4eZCjb5JkRA4pli9BkV7/9M7Pqb8EsQ5DI5+1Mqx6F8q9yV0+QGIjrOUd+SE
v/G80lvWlslIDtA/sPhwibYsst5KkUGNxc59nM++eonSkCfFVwP5EaVFdBieW9ul6Py39NkPIJwa
0tS02+Jj6IFoH7Qk7jQKmZnWw8/PKBZ2ORW7ugU8fvKjKgAYhRSY/vLI3eHUHTzErIEt/zTjPhur
rg7aW3GpDocgmtrmoGT6htmYLu03xUX2FqH2nzfuhKYBX6aBuX0/LpJoQcdvH/LBuvdIVf5BOCA7
gkHsiHao2p0BgaryZ27GYz1JPuPxl1tMD21HdKtKCI0v+FjP/3pXNja4KxaaSvKcEdNilxFEeSh2
WCg1QYa25r0nOn1xbMFh1rQ5ldvp8zGA/FK21zuJ9voi8xJJ5iRme4AVO7aKYLswA5NW7XXqAl+3
MMgebFW6Ofqz2n44zeu7P2kcvcVIFUmhZsWRsjjIWdJpGBuxRYktYi0GGb2kRfI4mpNKgSYsQqRR
tomVMgXrSub0m3OImKQX1BpTuXwwlchnnvO1YAq9mrJ0F4O/nxRb0UXL8I7iRT/sFnLYbpoRwlN1
nIbmpJGGbaifCXZp2vdEU404ysKTYd7lQyfsOGRzWmzv/pAr6M3iWnQ+5eSzF3BQ9oNthZEPMyLw
WCBonJj/3wwoD53NOaacF9fsawGVOuO7xsLT+6Z/7bKorSg4rjuf0Ixq+kciym6X3KMd+j99E0EZ
SbQgfEVfhpdxjJ7Qb5dcbZKNUbLO2b74uC8ijUdEqrwf+Mz5rlRefQr+7TW8OaOG6BwGJXNXRinZ
tI5/0wkvtqdgxi/vJKC9OiE6FgX1vSOlCSAK4TOI5NJblbDf7qiN2yj8kbE8yz50PHIaTTD9XTnd
K6GheFPsgHv8wss5YykskjdJP9lal2+D+bsSuyFlNM+ZimjMoa++zauNqzj+Gy8UhvEiPZdZQmbj
ktwKobjzp8I8d79mfYlGchogM37diO/WqxfV+etnu5CingMNwwrf/iG34WocItjy8I6bMzv0uEq9
YfSjTqulUH53Jb0ARgWUdI2Vy9bYkb5dS2IRe+Z4Kb4XeK43ZjhPLjRtMUfJsrSK2O6DbkbxiXDO
TnP1G+goKUYeHObOA8riGKnmq3k6DCXQpDxPamx8Sd7XkP3SsEkCVxKYIhaJgRLiEvViydaKbYS7
RqqKkRTMCEmtIEXDtWnHmiba/1BjkMRDilX7OoxqeAZczOFftx5tNVdUoGke6/+v96PaJOLWWefB
gtrow1BJ3PdYwnM0blOdQsJB21Y9rM6hj1CKaAFoNRmkGtTr+cC1UD693v/N0xDT7N/NY4UoRDj/
y4LoXw7h9r800uEGQJWVQ8YFedKNw6xp7Oqu1J6auyCC9cW4f7bbwpJsU3byqANIWyvUvWddfz7T
9hL1o3FnWJBaiMF6W9wUSmzt9GqwHJMw/+sTSaBPETgyXVJ1m6GaIEEXEGD9XTnM1RSAU+oLLMe7
TK9hTCGXbaXbXlt4tyBWpbzbatcSMcxwp9w8zUQ3tAXNib3G5KDrUJ3942b7ajWOo405ixCf3/q4
0XuDH21N6RP+Agxpqp6MZHeLPEWlFjvfZ+qsMw4Ra7Rj56bfayqu6Ibx+dkLDDgBXS8QBZedFSh/
ESZ4FMF6lYVML2QaN9i0tFFJ+9a8yJwk/E4yCRkyPMjpjfrMlT028kv9aKswHjUUKn3SjfyyjaWe
9z+I/klpnphH0GuaDvPLVFYhJK4MD4nZRB105FtwAdkHiUyxxSg9RWpl+Y+i9lBCpL5Uah/X648A
cmNBdQvGHDR2d1/TqZimqS8awGQ9xgF8N1R7fmhr29yNiyYGYkt8qLsdHnDsWM2oS71lq0fo1+zh
NU04e31cD6JIYiPKosqEOXZwEIi26Uk2RPTn2AD9qqZQuFf1YTKsixN8iYZ2G2AM3OpydPg3eEed
tq9Xql+ln0YAtviUAxtSGpELzEkWRLRiTyWZosZOueUMlE/NocSVrUz733DYn20TA8Jq/AINYFIQ
dvIhJgphXduv3vdpR+3F/LD69Q9KxVxLlswqP1sWOM3hg75ZHFtU/y1NsaPfTmYkhwWx0vZAEXCV
AJeGnO7aA4JK1TesSd8L9NXI5PZ+gMkx3wj0DEt7kGujkYUqO4xJHB5Iw+DYJBkpdKBOA+dVxVON
vmnw2U+/Q+quQ5UTkpctxITPXgC5qsaVGbsT5vnASzlFR2JYUisWxnv5HsmfTfeXsMwstRdbGRN9
q4s560Fx8C4nB0HJZkQ87ttrWav4HtCdYiv0J/Rh8e4mpbJD7934+4LT0g8e8Yi/KDLalioGQLuo
UA/ID/+7Eqzf2si0Px7qeAjYam34WPD2ZuspGd44jXcEqG8KzyOdJ9AcroRhnqRxSQkAFQVhl664
k/2Q+8f1m5QzdE7pAWra0nQhO0yzRckQ/v2yAbPxk5Gnfp02BAD+WrS/iIsQVuUQj25YPRxgfx3F
6jrfPfhYfwfStWJMiwm1yV4MfwM4xmtrNbdH4Chyj7oFtgVCRz7E9Q6f0GJ2lxhjEhZzW4zg/NRR
EnBcJHvDNPe8XC/xRuP7IVtaWegKT1zJg88CEg6wq7ioaCSx5SzDtzgC41pkzbF/D4dE7subl9mE
Z7YvTdKYnCRIuAk0RK/vT8dnZr5Kzvor4OA8kqom43Zvjt3xrXVI459WZjhxFWxpBJQ5fIqig5bz
DA44e770dDPdIW9ed/1tB8jml++N41Gulkfiu1s/aAr7KV+P5FRJRF1CqKhFtmmSM0YVDERLJjvf
n4c7MO8iju434ofE6lzRLJcNoZlRj4Axkx+FsLEuY0dg1O7jf/WYzLmVMFiteLzwPO03Tf5Kzz5W
noiWrsmgXA9Jo5kWAGswsdbxzCZ+aZ2ZEJV4XSmraWV3dGoF00BEGtSNeWU8Tl6+iruw9Xi6Tns2
3tvgx8/6jdact7x8TjxGjEtBT2ziNlzuTmmucSqcxve26TUu5WHbUkfY5MCcPrmtaXXyLolLWfu6
cXneYc4SVQwxJGn7LFPEtMqpAabcVIxqas+2QRPn2iIxRKEUQ7PNXJ4fNzXmbMCFKTTJa5eD46gW
Xlg1O0W6jxMIuxXrTwrlzObzOTZqdcOLiiO0TEYBcNt9YK0TL13tTuUMfzq9hzENFWx+nYq7CGpg
Szn7L+DXvnBAdywSocgCdcu/8k6j1mLR5TAAiLm8DE7kaVAvNZAL6898JRjzgNhdt4C4Ulz3w/lW
iEPvWtnGizuhufRXTjU97fMRRaUj4oVQ6JKZG6Hl7QwVRgifPpPRmdleYDjKVQwDWc0ffNpQrQ/P
BbFHat8ooIDDETUJ+O6FxbE7GjTM1tIIV6OOA7xgOF3ftiEd79KbR8auQipLLxdW1m37BCISNEY2
fAWeO8aoimMf3qu0QVD/Ozun54/wplIN0MjBZ8Fvq30AblWr6D/fsce1uL0jKyOy1meUSbgg6KUp
qRrREMAYAQM2wgPBD/J9PNe79zAUUORjNpC92mfGE6N+zYC2feluQmHQe2ICTaR8aTtTGzOuvvhz
pODejKfk9dYEjWwPOHyCB66aQAbat1bz/1e5l3ChmyuVshnfoHZl1lIjQ5vav2WPvQxuynpCmY7u
PRwYZDtmqdD/R9L6XO076DLsMWfEq277P+DJCu95eUi0jJHkRL/ipP49t0ZPppK+i+y2V4T3kxHj
MNgX18kU5EsEdkKqSrf8S2rIXHake6pTPrICRdO5QxwAoKtr8iMLfNvYI243tYRrY/QHz5+tO+gG
0w/7NPf5xRYv/EuJ0ZyLbvehsDpsj38NsnM5i9CnOLq2pRHo69rsxooB7gPUGZCh+9MT8foNGJqi
l4InHalIFMJKP5WH+2C3GKQGS5CsTpb7YtvnHVq9GWFQtBAHxdFEyFooSwCXeENu3/VGr6urmnKg
KaE29ZaVhGYjwBoBSiI2z6kaLnFcvzijXcmOA980z3gqquyg2FYUCQwM49NYPvRuIFdx87TlhbYL
JmXM6m3p9L5gzwlEZZZSx5Hlk7Xze+9+uAuDPeClSPd7AodArvaTk7fBeg/VEbIgOFqpubJkZ9ao
COnXLEngwBTg2yqJ29J6GIemgk9kf1YJRCDIknBU4wTKreeyNSJDPecbNlJ/caLloqewJBIJXzSJ
Hoz5TcYdSbmEkt613WXVb/hd/e3MfV94C6W7iRka/htQ8ZuRcHkMp477o25+/9wUNxxwJ+2TkOv0
lb0IVEW/zcggENk1r2Isy3YVxMv8N2owFZ9baUs0rL7STwohT6GfHsZailtr0ba8xrQzoHuax+2f
4qEgp9NdWBVR3+jT7NCeynKuvt0eZ7buKgrZ5Dlg3MiKc434qPFNiX+2iEz3D38LlMdh9NAPaepu
4EcswbWBu1xP1Rl0LTXNzecbuf5k8DyC4ioS3MTrq+gey3pJXabJ5MtZhruXNdhxxDzSwMsLODVy
W46fCd7BYKj4ecR15twvNfseOSuzySQVWp9OeA5rx2dqWvXOUT4LYXJeyEGtLQQd5Iy/CKwmljMd
1urAmt0NaCEn4lXUhxGvW2jcPK90Kmy2IkX36yZBneaEEdRJiKXedZoZayX8E3sTnHtHltz/bzy8
v+5il35Grt6r+mSO3w1D3uplAagcNVFfW60huPS5xN0q95zpzhNBdYEtMCNdO8ixpl/ZjH2tubtI
Zb460GK8HHU1dSwHg9OsZZYI054p23EJu4NpieWubRpk2cYOKof8JwxftFnF3H5AJxjh8dFC6jUf
uijEaJPscUMF4pYm2g3qOTrSroXnGDPveJwwbLI74oS4ZpvtqgQjBycwMXO7SkZjVXRooXHchsMl
xWY/0I8sXQrmpm2/4qnnKi4H2+prLtQDSJrevI6sUh4eil2jc+C9LqfybDstQmep4MZ1HlNKMjSq
JZWdPe5jY5W1EwHo6PvzTS8RguWOHnAmcomsYBtRpATmhyQYuZEEAS1T5+ErggPEOtESSORG9o8F
OJ0Mn9kfZHHu+OnIcl6lMEcEYRIpvBQvV1854jZsNNhbO50gGWtvTGEAljISkCAHlcgyNHFM31g7
txzRFfwARVH8veSiPwya+B5W7j0aBi2a0ZxJw+hO1K/3Oysj/HTo/ilwd03XRVmXqWsntGM5aMF5
+xUwpotzhsi/9jYomveLmVbgPJ+0YI9HsSDfKFI2EUhqnFRcddGxZGiAWBWzu3TNK4sXk+zZROQB
ts3hG9GyzE2ru3q2MYtk5Mw+dlCZCVP73fIt/4yZAa1f7K+9Vi+sg7ZpVP5x9BaE15sK/m0Dr35u
S9+hMOMzN5+Uzo8YwI05B9pKusMi0Sh8iq3OtNs7lS6UZAm2ZPMouB7YSeL1MIHl4502YampSIv/
IpxeAZw/Kt70+Tw79okBSj0BI/YdWNyvyqaYo827xg9zxgTr/etO5Wqu6b5UEczOXH0ZEvF6UjUx
VCE0H72s5y/+FdJWyPM5IZjIGXX34VKvIZeRfhktCXPMJFpztibp2gMabFs55tkdRJWb0X0g4HoY
sEWPrzzQRgvFD3jOu35GBPcJs+OdFV5M7tx91S8CH6oWplIGJ6g+idnUCV9tjnNwGq3mbwMx36w6
2UhHeCJ6H9NPnw9narM3iRf1KyYRyTWUPEESPEi+jdLv8EbG3XadzpiBd2DzdE/y/C4vFTc6lnso
m5FuQS3/+OPBl7A3P1R7YcslvOs4opuNBG3SsaMZLWAl2Ff1V50JpVi6xnAon8wnwJbFG2nuF+eL
Lx6LGM0i1mllMF/8oJe/13/Pkno3PxUVJmka7VWJG3zuBhD8/CuSVDocXFtSHZyv8LxWK3rwyoK1
iGVbCiWiGPgGMirsJl3QKSsAqydMWXa+fNGkHiDjEfwJyMuQ9QKVy1h+wIvUpLdy726QLluSr/5V
OmnT8h6waI77fSqCBECnexfV5XGayxIR0WPmMNgu1fzevq7UQMOYiD5OS47Tp8b84w/yjLxRGrKA
qjDdTbKsejz8iI56viKLHUzREgfMPC3uELLJHSgPe+bZInNErUFlwlOa3IXm1DNP3f7GKmgmG1ly
To0QULWaN50y8eyuzs0i4I9goIS8KedDnZuzMrkzvvD8HkE+/VCQhHu6bmvfke0jbfn7Y3HcUEyp
pUA5rweF/fsXFY1flYNM0lnNywyer7CH5p9t7NRlTm0aIO3bkRFpMj0/MEm096UGpI9CJuxsrc6U
H4XjIZY0fD7a9NHyl/bkbJoODY5344ybmH7jcIJV9yGR/+1OFfeX8xBXBZdZy59dxe9U56npOUe+
hrZNNZMspGtIWG7TuQQ8YIfjGPpznYPjFvPbS+fgR15T92oYM7htTmpEJdKigkFnzXmMEF13kHoP
jLVXzxmdoiHNaSLEqAMNqi1ZTc4HBMI5dpMd1ZeHNO3BE25A3bVct+V2YGto5CFjchiJwtOBX3W+
t9pQ1MZ7nOtWfmF1Y8HHlxTk/rR/syZWNmiOeXOoglZuPGuzvB6gHusS92fJ44q5VjqSb82UP/k9
XB8dKRuW3lMwMpZWSbSgvxDJexv9Ua10gzliKBXymZdhFICDXwWYiaMZkBC7Ic1vpyK1OQ0v6XDg
VFiPB7pS/vq55maQXTSVrXZR8HHepR2jbRcA7TaBolBN6gu81pgDgwF+CCCiH2U5nOkPVonwaOF/
O60oEY0uqEVO22rCrulM2gNUdMqJNC7FFFvSSbt7sHpIMV8jOcsDzpmd/RIuYglhyaE+PVh9+eBs
JRIQgVE2l1aE8aibMwa/pDcsYVvbWM3UxX3uQaJWFytDCUV5gXK257gJYqLRl3as2k3NpgPVElfC
5VKTNWn3MgyxKshIDHVyh+kVBR/tNkth+RkSoPaqCBIqcyGAinzQJU8lcd1Yt78DJvy44Q5RZycA
WzcJsNJXkXZ/6cpTvOJ98zkLCzdXxubpYHPauoV/s/CD8z7NN62F08UtQTlJqWZybr6wLthDCLE/
If4ixyCYYHuVPxGkL/56inpwYYAk9PbVRHFnukRoHqCmrYwc6yz/dnFH5vQ4bgubKsCzqPTinjY2
Mh8lzfQUBfB6V78XGj5sAJmtRT0dKLcHqdy74dh3VzzNxD0O5tPS7+vXeGfF7Kw5ge2Qgzx1YPAT
nYugpI3OBDHSZIvMImSapVJH+fBxzHmwQSWac1GlLm028JUszBQ1uG2iJbl8kZlZPpycH+6F+snh
+wQRKFrQwdIDy48InSLLsTWYGWCtsJcTn6KS/5l6aP1sgHaJ3VF3FQy12Ldo/Cv0FrJD9b7HU6QE
Sawri4leIXoZfd/BfT8IV+USzdyghknC7jLdiMV009BlKB2w+404ZnLBXyB+vmQuLXOJfxsXwpxr
o9RJ/vYaSxVSZq9R+M0wh6dziMfo1ZuhEfABxRgSQUbDpb0gPeg34/yQg65o2EO+mttum5JUPYtb
lu2mgLeubr7jITkDv5QLGmONBDRdhAHh/64jICG69QKqf/ueTjWzam9ou03eI/oAGLvJsrWvV6xF
uC0w84/IMHwmCDYqapm0EwkMXrh/zEEhxwdKOA6QNevNbtqOozO41UR5cWHTFs3wk836v7bL19Pm
TzSI2nk//LJfGwk7+sWUriRzQ7dBJGSoHE8xpb9NlnaJzyBVllVZQrVQjD1R3jrV5R/gdvp1osJD
7vI6WRPcOQWgCYhSKElIILAnHyWrrveSxR0oCv35+NX9RWrYbYNlcT7yI8uo+I7zt1T2D8BOrzNR
RdLuhRi+waMpuABgkxRBQkAViUuxsO0OG/TYJStcGXEUkCnakQy5FSl4mYIR6KQunr540ItIjNJn
e9g8hBPzXNrvM2vQ9aDodWkWA0YTnadxA/zPKYh5+4s0X6y/cSO+KzQZZwjdcuwbN+Y/VBKm+Kix
bjEhp2/Qj0k2txP/X8BPuGXg/amckROu5BBV5GA99NgJ1UNIiOYaCoWuG7+dzj6XT1c2cn0qQQch
AaS0j53xaHJ1V22VA2Ha88EqKS2Gc5C19yVIRY0J3+8GOY/eGY+T9ZPZx3bHs7MtZmZVfQZVdvap
pgulfC/MRC690vJSaOBROT6vzZRjKMatBayqbtwu0o3hbQDx0vo3ow4n7RWi/+sO8wc3ZyZmR1U4
7FPDmaaxgNYW755cJVgCok6tJ8KjPkf1XBrBAvXpGT7sDVDAaQj4yMBxm/0u8DEafIcJWmbg26Z9
nzl9Z+JYyLC4HVlZGoVtYARyJjs9IoP7ZW37jVAg//kveqp1WU9proeQ7EM1JrcFI7kYCDZZjk6H
op9+F4mM/kvjTh//Ud0oUvVWydR5XKZw2cbA5cU5SqeNjDvnfqQFluFTNK9uSSGzFtpTU0GL8krF
CJWR3uHIsl0tTT5DRMY0+pFzbwWWOBZMR2h1vS3KxkbQOT52jWXpxdw3uywNRd8jWUdf9soFSZdF
+IlzvaCTXDzHEtsQy81oyjTRNmYrvwqyjn4GbV8oG7aARJaFESMCmLIJE1r3X9r1wVtJtFBWYVub
MGWyWdLfmzjAukFeNfGxN/YoWnVM34ha5atWDh/2rpyR19W3cFhO9knl8/mnctiy3X0vn2piMVP4
zvE+BEJPNAK5cBlhPq7Mvm9qfwEL2R/8rc7h2yTXGVtwIoSXr/xhrTWB+JQF9//7Ck8bqLr35g+q
6GODJQIcdRW7lletPX4rGxMqTRNkNhTa1zzCDLtxIoJE91Ha4NOpSJ4rWlldWXKHKtLydN4PWu4y
JKrcmdzcLXZhFxdNK9jV0Meg9NWDaXqHGR3qEwiXusdAfScUYm6fbvCY1hGxuAdl2gB1vFD8plsC
O07jIBUHQnL54j06Gc5xjazz/UOV5jYmiixm9ZLPE7dPYsVynvIK/h3id4cV/7Yqp19GPkpZ5kvS
t/f5+z0Bhmynp7f5GOfvkJ+IkeOMVwQ5Am/YElwDY7yqhyCMTbJzv3yYGpxUMJ3WcrhgvLG1wnyC
7NzSTLwh8mM3s5j7I/t2id4/cFKvF5v8lDP9/IL/fOHz07cn4mUeW4Rdb37NXVtGfIufduWVi6si
5PABv9ltolQ1d8wKx5teKErRPCNEhmjIoIxdPRBppp4+pcPh1uDfrP9xr/FY+OHQxizjmITc3S76
B0lw4xweueed/PdAVHMC5y1fSVlFE0fpm0ZgjRE9IltFWfAaSFuDWVDSc9UxBp1jU+uMi+1ABRMi
RySgKVQbitValEYX8Hif0KXwEiiEA/FcNB6uovuWE7PGAeCENL774deh8e1X2mLlS+lhbdqWQOUj
/amR9raBP/wmdqezMzseH7VE/t/xtQUOvs/++8b2CXCOck6HCqmSHihVE8hJNXxk6ttU9gvNFnye
lBzvHE2i3Ow8+VQzSmKq6cXCe7P+4mRiv+56FS1ivinyFGEKDJop6CIMyka9NLnD7Q1AyQQJBTqi
gELits7pVfyevM1iHdQlK5kMYdTkefR4bY9XfihFbQbxZez+XC5sPb4YcXWjD/B+/u3oIfySCdmf
ZszYPymzL04FJJ13wv4rEE8SAvJZAih3oqlfCld+rFh3EUDvtzKNPo4pQGvYpNovT+YqsIh0UDBT
Y9xMsI2GvMgunW39k0SE0ivTkZcE8bWPvECFz1TunKFCZd3Vqphf4jyu/ZgRYxuimVGO6dDIy5GQ
9t8oNKP61LgxgtHa1Uve0XzuIOtknvTkDL+h941sJZELG7vthc/3EOxwHGcJG/q0zVvqyEq9yZ/f
o1XcSyK8Q2q+ea4dRBouwpji55yq3TKP/xcS7hJ34dp5d3/KE0d/+RrV6esdetz9EMWDxutLLMpU
8kAJ7Lq2t5ubHA+iwCUjO/bbwnf0Yk25nMo33JDpnh0PGxpYEMYeHZOFzjdcgmEMBugKBakPZVZP
zc9cjdUzW5IHm3tfHZbzGZxTu8bx2lJE53RDp75ABbMn+QBmQkCouJXVUQ4p03jrwh09xAZ2VMpw
58a3XKoodWljo84xN43gBjbvXb0m1sGLANHPXBwe6V6bKBASJx6IVkea2FTiEdsNSI+NeKoP4xvx
nHAUBdJfXSMxsRekuSJEQDYWD548adz3m3J4l0JaM6xS20fjw0o0hR8bojGuzjrn8s4tpQRefdXf
jYzSz3lccGeJ1KN5n+6xMW9TF0PfoGJb9QdAtV52iDx87vhWrhpXePPwbyUrV3uhAbX8gWwkRNyr
Du/sUxgEJA4rYZqw33XnEVjGa6Z2iVqFc7+LjBSsc3QExcgEsPn/JgTFS5SIJQTZh3kTPPlyw8bs
78sdbSwVC4ukhL1lrF49stSMn2UBGDB4+8qW8dLRTTCn+Ra7duEYhFcQYvnEPbB8pEcCXQYKx339
yIL4eDxQwpDQVnX7eElAbzAFOqRk84NohmPF9edZcr0MtqW/NKMvsR4kpa89lTK9fPlRRarKl3kR
UjMZ7geQ9/6TdEo6126ODEjkNO7/JusPd+Jy3X8aoBEH77swX+61YjprxWhei+NWsgoBXihGQPe0
wV83xO/gTZNsoChdGSVkbdi/9BNsbqKycWpfZ/3V55MPUZHrjDXIF29Js1LFuVpeKQe+B2JDmgl4
A+3oOPWbm/fmkE27Oi4BfQ4LA2JKTwfLCyFxE9n10cTky5vf86Zp01+y1AFGHlExUkcn5jLe99MR
RYvxs+6FvMiSERADhuXGfJ0zQ8/tsWbm/WfpolGGLKeZwyyIWbxAd5D1XneKouC7/gf9s7UxDxwJ
JW5DcClCDnXDAUvmWVS9vCgpAsAkTXkTc5YG/31luUWE7cCeAoCvKxP2IhE1O/O9+a2CXaGMOQbH
bz4u+wOhTNwSuZs1Z/5K1sKvUHAC+Kk0+KYj5VpAT+HtN0GT1Tti0XGz77Pv0APdHVFIEiNZpoKD
YznzbQL9xp0lJT5wNlY/zn0BT+ajLmB/zFkKdU6I0xZDcu/DMgg0wAJ+Krl7GQ5ui/Rbiu+yxV7g
+VQQPwMc+7jQuwxW6EBSct/vAwiJZmOBoTsr7bmRay0+U6uKkvFoHwSMYtOYjRk4Tv1LDENq1bey
68IigmzxCHer38uZar9254vc6s+Wtx+40xXbcm0XwoddHXpRy2mF3ubAze8K3JxdgiFZ7J7odTdQ
x9x+x4qoSMamXAYRdZ3+UM1z2TsrIhaU4ixZhEqRrGNX2SQ4k43Jh1C5kP4fchaseZvLpces9dLV
IuoJCQUJ7FkMlZfW1blqyFxBDSw0zF0IqD4QloLTCvfzgAgdSBs2geyYfWf2cqPZabJO09+ogJOf
8s0St5RufDFbUTAo6L1RKRSP4kzVLwIVKYyp8YWVb0cwdVPQq62BmPzq69X9bQ4rsr92lOepYpHy
9+SKmFJIFLoen4Sqc3ojoGXa0/vYQZOlSySUY3QQeHWwT8JRHx/tQ1cchQgodN8Bp/Jr5rZWuXfW
QiLjUI3TnjQ/9KirCjotuH2LW17Iou7U4HV6H5avw8jeNYp9EgFkZOvBbyp7l/hPP1CvHnMw7m5i
BqTKyN17rc1wFQRRMsSvqDI77H4Vay4NmWcVPENcTUSdXTYQCmGAr2XQ+GBaDbBg710OYjVrNMLb
2rtAbyn9DCuBAqb+1jqglXdujtrC7tOyuxWk67NSu9sQbXS4AEG5S3yGUojCIRcOT3L1klQfEOdu
6XeN1+aZwPVqVHkNXC8qbxk9tNPlWub2nrXUOszdD6KoTFQjbC4ZaMZ9POAxfRaJCshPf9C3zqXf
Ex0f/Ir7ylAJ/00LKJztlMfL7h4R/GN+y6CLC2Umjjgvflc8Z0qCMQQO2XUrTDWvC85gUxRRR8so
f3GJ6iCakVRusI0cISQoKmYh9hidmFywiemPRFGawFa8gxVGlUM18iscNI1R9GDjgSwWbxls/i0C
XftvB/M1EVz6djCP3cwoB5tsqqTnhTMSfAnHknNkQA9TzxbUFRhlb7uR3M7k9Jw9CxvRhr54ey0+
6nTaaw7L3bZK6wwrUSgRTl1kiIDuZZ854BKAfSgoYkVm3yxGSrLCHU4i/Vp/+aMydNUrrE5aoywO
i02FS7kjjtr63SCAKsHM3dQ6zt/tHPajE4qQu3O9WGV8l1U4etVNQk1pZGWfKCbk5sUdrHIG//RY
njvgjg4ua2xLTykW41hkQ8lBTa3uJ8EcGMQQij8tBx/kPpuFSaehnUYYtin2Aczw1DL+bOltHaMF
QTypUO0PqfNBH5KildSdjZlsbk4sNCYky77IjeaRpRe3OG47mWOIAAfOAYaWKrr2f8WPI2sfoGbT
Au0Qs7RNT8OEL8pnDilenaNuWW3zTT21Oa/2jH+/MBUr2494YeI5NJmJIsggo/FppicIKo63u3Nk
BGdpUsQbpKUq1hmlNB2DpuOKi8rvuH4m8prm3IVUuBdO0MI9ejjmPP+0waNRcoOtTSJaTrbL90SN
gr0hTL/t2+Rs1nUnJzYStTC7Ptnt4rprIVMKehfhnybruEBLXSCzPOD3sX8P0aG7MJQ1Rp+4wY7s
39vPaLax4/Lfl8WUPD3yKNIQfmEEYxMRhDKC7wYL6Bzoryb5H/42h+Kmqq8IHTu1LNxGENsru2wC
BCWkIyxyO45hHU3R146gaWi6FZxHaQF2ZoDZ7YusthpiGjQGtmz3qcnNCBlh7bLWLClXlCuVxHuR
IGITVQrQ6q/sT9u90eGTAPNgQcJHQm9LuMf7DyEQ54a8wih7mRLujnMnoEIEPrbAvAm7kPtIDO5r
5rucNnvqLYK0ikusKwRjl4aSAktOTRQG/0YqcV0/WuKA9VG+8s1ARFvLnsLvSUoySXwuFtqH+AXu
pjz/Z6krH/qqNCVqncHq0/fj8wQxCbCIJiqSXXktViOXTG8FGupQa0/1Zkcsk/NcTm9YrNI4qTUx
1WOIBAPn3zeYCVtH8EnvrQw4CylkbYn+Kq8sgqFOcrDUi01PcTdUf5FYIKVqN3oXIJRMuMhmtjYf
6cbJgQEA/+mvt/LOqzaG246VDE9HCV3kS/Jx44PngROO3ltf16z7AWbfjl7ufLkWOOtIPQb+Oizb
o0fG67AVWzOnvZ4CQAk7NBg3/mXSzphFCEy0RTytn72TeZjuxAPqv03CF3ptth9WMLfR0ZXuHecn
XJN0iAQfucLkTGTkRtRHJizlhyUF9jMm02QAVSvUFgrd+3bQ5mIgg+3f8yHx+gcU++QFvp/T63Xh
1x9ybrIFvN8Xbk6EJKbU7VTQA8SAXtgvZaKSRZi6LDciByzMAD9PFwYzEEQ0vlmGiZWQjysN6Nxy
AfitHDwSuoXqY5qCbW8iH9NtSIkbrjuvhq1f0PqEvyb9kyR3nhqkRFVjWTDNwxWwpgOd6MJksF6v
xQiF4XdiRD8Of23VMyiynd3r/7LXVZ9ASqNdtitF/OjhFW53Rx3Ovp7ZoaoWHUnJf4mC7bud1XdB
0dugEHZKVrfTKgRBgdfcN9gmvwFknxpcMMRiidlgUKbfX0725mmi4capjSZuWcDWKjceEhoqrZY8
GmJ/9400GIaGICe6BbnuQoKeZvNiyjMM3cacB0uB5K9j5kyMzACLs5WMhIHezB9yTq3QogK5Wg9e
kF6E9A3KQgbsRl4lBbtGXgUgh2VY+QbXPZGare1Lx25fdX3ppxGKCFHJM7irdpXOuMlAkbDvqz99
fhyaXLUGoLuPrkG0c21uHAdocBySSSZLa2Hi1bjV23Mj6KUZwAGpqcUwcS+s93YaIKvnaVnV0ZBH
6vZMNjVy36zxkyDJ5uv7PJ+/eigJEZ+waBE6/wmEvry8cT8lSb4qO2c4SHs7l2i+aZ4DF07oSvUD
3XyO8lA4Yk1x3KR3cYDCZRSYJKaFG/YKFVU0YLyc+rTHuvk1Z4wQ9YpWWCPOE9132q2y/1Od5Le1
wu8igAMlwbiFQEY3BlnCJd8D2mm950Q8t2Zi1CIpCDZimtXJA+eJYliPw0eVmzX//cXd6cr+VeXD
6ZbDlbW7ij5AxNDoDV5wLPuGhst7VJG8P3dEbQpIM1PORFM19s5w77At8ProVM7UKPg0xjCIBgYB
CMJWduDCTgzBnzJy8nmWCdOnDhTlwkoWjusSNif4sZQcaF9epVPcq8ZY6+iZ5waEP2szApBogYWf
lWJs9W4BGFj5xXwbVma8dLIWB0894o81y9Nvx/6GO1jaTxM9KjuoEuuBcdEOmkD7/G3TapExFQYT
x9l3YKp5jryHKjEVmiWgFJZt4UMaqhBUnDLBNioijS+iAVPZ4gSJK9zJAaPCUdFGVklXT4J442P/
87LZ9hxi5//dkjFFn3xAwJGNimVNHz60n3/uAN94OQRURhzFi9mtGC2AakDNyxmotla9jICESGw5
ZVreUaIbX8aD+vUILD3WQmMXCi23jbAm5mb8mA1Rh92G0tHE9C1uBy/tk997vpLKpO2f3lFB8uLo
H85KD/0a+j4/YJtxYBNKgUsULp5j//0JELjN+D+AH5GfJ88w0vsZoW2D1sl2ntiB62NnuO1orT10
XI/GlugYn3MrbUyb6IiYN8Y+Wh32yvdEYLG9ZQ0oXwgc2XgvG8mKdMywIgPP36rCVAfnjWBGVu4c
rslGCbD3chVy84v/LO79+xXpKFRSTvJelGF4dyNSZfa344NlTGhOJNKqMUNBnJsXpxTN6Iu9COkf
1JJO2JeYZU1oLCFSLrYXv1sFdT3bqGKA3cnLN65FdaXvjJ/lF2k68Izfr1ot5uhXDiRhFeUSQ7B9
PnFVAh0qPH3FQi1+L3GPyERPR98JjkLSzmrYee32nIiPLmte2S1TxMDXZN2mTGjBMvRm9q1C/uOU
lnB0tDuCG9PwWOwze8SCLQR2bFiSi08f41P3EdMwR6+c0ysw2e9jIGTqXU83nj7oPyDIvUfdWH8n
0bTHUxrv8NqpaurUl8+ZaldLVZ9Z9luxyuSxerupuR/jHu+sYaEh4F8Nhup1KkrsAMnUd3q4ClTg
8Blj2DWfvAraygIdNFS80YOebnc+0dp+DkhBoelgbZzSyyiAoTAo4WFCkWr3j42IXjXNGxUQ7auW
mzbDPO4diHHEXY1+hrkMfyZLPrMkpWpMvBL49gnRUHR5GW3+0BexXPTuecynE9WPsqlYe7i9etLi
p3B0pkpNJnbdS+AC5ukqfX3wv9HuTmaZ3LhcBOMULkb0wnL9Ya3/Sun7wf4IuHsFJHtBHhslqzkB
0NMxFWl30RCcQIB7tLzNczdGaT+TGcnEp6UXjc1aXyvl1YQzQfh6XI7dVDOE856I4sBMIqcjHvSU
se3oMaUz5+FC9Km/x8JPgJYAAF3qT/aG3qNUc7FW993nTARZKycjT7uGqw9GPUfvhJ1QhntCcypg
uAYV0ZdvB0u5FV1l6Hq1km5KhEibF8rsyu+/cPv5xFP7YKJZNX2kLthAP76qlQaMjileZ2CwD01k
NN/vZ+4KhC2MbjPpLKJm2HB0AapptL80ZHr5jEroMTYYGn5Nga3ZeUkE1gw0+h0DuSIRxB3o3T+S
MVLI3tp4O+KbsgidDFXhGF/33UZvJWpyYrHM9vEnn1V16lRJ6Nk5JnmdliPhG1seReXGHm9UsVad
4zzVePoYbSOe4lHz72xZhmnLJ4uLElP516KKIZ/ZAsuqQH5UHyHpQUN0Pb/ykWzyqjSBZMC2FAW2
PzYeNnTCY9uCaff84LJTvilj7t5A9AHCAKy+mT0PZCuMDh50AQUomulWEhf49xu3WaupGh62E9kn
omQRtwviioUEx+fmgeg4AYcQFHKpZvkKp/6pDCE/Wt1fuBfW7/nnYrzWdOa8kmdvb8gdrWlXsyhK
OohdmmN8QvWLwzDd8//+wMPLlRdIUCL3SqEG6RWq504pLU5FM6/9FyWIuC9lvG1ksbENP6DzD8wz
zz7Mz8mjHnPukdeGlpXNyo9NVzZc1eDPpdpkJq9lz+8hxo+I3w7MOKa7lUHEBFhy0ZEnOLCN4hXM
PpknbsHyn0hLBMhM3RlyiwCh+CzOZEvAvxsIDtKKsnLS0YrJzOWtbfawDFUk3c4/aZfJRGzMX/J1
wWVUY7zA5KQVurnbi9hUbBl91dPyLOFIOLa+q8UeM9JO4tUmTnixDQ+Y9x3DzvFWRth6cgoAQ682
zdXCq6mgtAaaDbv6Xht6I7IL3WmFuPxsTx3sfAbkiRPmNrOrPRhTjTOortBrHTuJ+kiG/qZOGXtM
x2MfSwDTUH4rBUmsG8sAVSjDVQFxAGqgsxkzNcNjdVYPUfwYvWk/k0uhJDaVDaSCS0GP9oUkOcCU
oPY2E5Lib0BToyCOBibi3QNeMALfUd4rMc+jSC85We/UMssGJO05T/G31M5OLWYQWD7JyopjX+eC
hi2AYz5QW2MQd9mNngm+CuByGagHNaUTNj+MIGThh3ddRBitfTTyLp9aCJGHjrDge9gl3vCkZVPg
daS1d4NBrA0szqnQWXYZ7ZdLj2eflexjJy/tKukUVorNEMGsdzpvYRGl5zz3AxTCa3mSVXiORW7y
pCY4sKNnUzb1BQoe5F76sUUZ+a5cYUjfDfS0KNx3G3+NKJRc0tLMRi84h4ERdtdwzh2HIY8cwFbz
mU1/liihL4xnr+nGKEWRe2FjRj6YosIsFvXJwgcuU3Udy0tw3ln3o192F8ZuhU9dMrW0s4dwtwAp
13c3jnN035T9EuiI4n3MpmP1NXQaYK7z3Xg49qjWnfGKyHTCpbgyVzFf8meKYJbehsmV7eGyTnXH
7BTpl41GhS18k2auNL8PXCU4PJ01LhkSijlXPgC8AVO7ZJYCK+3BVpX+RIg7OD2KyAQ/ghvf7NP4
2CQAV10DKdsPzP9GvoQv1099eEmDxZBHc1HmbDvQeoTADIRiBVPhXlz7CM8wqJTHfBKYixsh9O8q
Jwtua/hcrkYytjIdG0y5t0/EIxU1EPn7qDQljR1JLqJBm/D1ZP9zcchmsf1X1JYV0IL8s6mMP+Yu
9VjBSPOTliW+ljlDR7J9EdbP6BXBXE+3aeqYbUM0ROpcO9Yh4hT+m3Cao2yEZmkLJi8327icRXPw
OmRUrhA76XJMucP4v+ZSg3s+Ci+WuJSlJ4Sd8e2H78QoLJ/QfJTXcJZuFNS20DQNErO3Vc4Lk8xU
B8e/uoWYpZgQehqOMOiajzl3A9q0pZtcT2ibdpOu/+OGAL4X5EForpdInpAiYWYfDrOmQDyB0ilO
yS/OzmubECGslYM/UHhSki2W08HQFivF3L2WcG9YlOw7hdPnr1FIrcwbvGlRLene2i8KScfwG/ny
/RZuklyaS1aKOZBi9A/Mo3GfRakaY1oJ/koWS3EWARc6FQzfMyzTTQh6KPxWKqFqY5SOf5obJawV
O2JpXVECtHH0FMzjLexM5ffYHNENgAsl6U3G69OoOxOsvJ43I3ucqqPYJ3hkR62jOO9nh8288qBh
bq64O38Wi5BO/I4A78hsbq4rAYexLvLzAU4YsRs7Ii+iAGicouTP8vOh3xKisiOqirm+RswYXwiC
03HPoxQ6/HO8PkfSqyFJap7Kpd3423m4PpK/sn4U24C3FpF+pTMPYSlq7SAIZ22Yc6tjPv6z5g8p
c20fxtuwttgV++SmxenAKXHcUORnbhLyObTqRD+KWXStGNv1vvrkZjQBvlz4Enzw2ZStm3wJPhFk
HLam6pFZMlv9iQgs/tLKiRD7BcwFOFL/AJtOcoVuSTgBP7D9y9RL2TLkEtCKYDZxMHcrAzhgujoD
8h3CQrSEQ2cDd5FqZEwGet3HlYa0d1s0Bp2zogPLbI5doZcT6dsRAeHCtkb8xKAXp3glbbnQkau1
9V3Hxlb/CjgGq60ZTcjNWxRk3Mf4yfDRlZRaNjSjgX6/i9/XTRit4i2+nKw8k/gZv80yBFYSmysN
WSByTyxO3Vmbt2wAPF4x+pEqTnnew0j/aUKvRXop1b6Rtk5VZ47FULbI7YadPDvVh8Kwiy78kkxW
2e5MrEyr2HS7RzY6PWP7/mBNFKbjVzeVZ1ghb7puJUMYBppnXaRv+4j4SRu/002OPXiaWoKlDsgf
KsmPzaWIKYb06Q5jM32wA+/EkqldOt+359uBbBFA4VnyUVBQ5UKJJBGgkDppe47Bn0cBXQPFI90A
acL4qARhJwj/wS+WW8FMTxM9gcj1QU/jf022SoHeTYzw+JovZwuLhmGfFdDs1fiJisVDjMsz8p8d
D9UIVXWQKq4xByUST/YvnYHyNlPTS+sDUMOERf7Amz9tPTW5vBmGSQ5oXy9fpULv8/cjJgBoHKBh
QCTUzv3q+XaMQVXILEaGe0BcfGfkdMr724RhDkvajxgPRXkI0mRA4qJh0tlYASlWvg4WxDkuB1Rv
nIOIGg40XHyRnZsTUU9L3Z1tY2Eb3RCM277/O+IMMWRpKMBDbR9gKZXTUM+0pBVapflLAWIf88/w
h/tEq2U+s+Ldo7LsSbwNcbcm4a5EoIhBp06g5a8iydWGcMYlDAID+vZMsBhXg2EjB2Fn2TWXWmeW
NZW9dX7B1JG4l9p7Y0CAlG0wPLCwZgDX7NazF1LIdBhCsiUDjQ01fBSe5kLtQz7kaFhvHk9cch7s
LPKW0olwp5C2zy2HH1lzCW+NhgiyJxVlXK595u1hXX3WPt4eh4jVAD/AKfbHGwMUErCJo+E1X+1I
vCIKxhzwG39CWxbGf6LgPrDegK9vgz962eT4GMge6oXJkfZgNN3Gc0lJHXh0l05OlJ2uEBfoU47U
zihTbSgFRELc0OfVVHVI6I58WtF21x/9VZCjLIZjd1ANAzSHxf7r3aqyZACWa6j9yOPDyTseWfSN
UzHExWNWF9Czg7ZCwrBUQ6rld0pQ+qYkCRreWOHAQeYbRjC9IeOqVF9+yLmzaxgxZa8qd+LlRM8j
j81D5CQtRCR4L2ZGYiG3s9qbDWRKLngQezeGgEhLp3A5SA++0KfN5CBhqnew69fVqoAGefNNck1V
kbE3ytDBuCpphy3sLui0Fe0Tvgi0Y1N9snPZF3s8v/R+QXwXit4n6QhPCYL59WP3toEgXj0StzHX
YvYZx1Vkxi66KpzsX19/nO3f9f88RHY9N5E1cvBrViID8qB0YGlByS6//PNoFx3TiwCJIpDImXZ/
fqJcd2teCYSCcVF40U+ag9dteQ9KvR/eQEybyvy4/MbAJEGMlJbSY/conscaFemQymvTQPCcX3tx
XwuL1+Vf7lnlT3fT2VATKovTAQz+4F/gHRGFqrEZN8/EnWdKCSebgRrh9wi5qYY6ZGewowjU8Nma
nCFKCOwU/1HyHXFFzd1HtzmKk1BbQtLwU4wVX8Z+M1GsvyejT4qk97Zyy6VeZvNaHHkuWpOwELlq
n8To3quMLdk2gXZTeFoodhxNNA1TICdBQ8DHy5/9QPolNFF9wcfFbDWmnoThDlD/9xljxAugKGyA
X6yA4Y712Ne26+sxM+l3iI1mVhVPeGLwpBDsQ02L40C0eaKqRrzeaLQ3ClKkzGCeuUSdbOxgV8J5
6rMUu+fqHHRsMYSZOTk7fsQkGIBc79jw+FBomnf4iXHQp6aBqeRclzrWjfmduA82aJ1bVEl0ob6A
xhYYbWC90Mqmk3Ct1XlBhqkZ0gHasydp5No/FDQz/YGWF6XKsrKcQMuCLIM/Qh9ITA9qGW0voZBK
YdmYzIkG9rg64Dej8y9CGVLaOl5hksQdQNLeTQOL4mdg7lE19sqCFtt5TjRDAiqkT9UkZrWHfdl3
AL0cCSvhKqxSR4jygyOkABVPyNySKtO8YlUE81jTOcjQeyJP7PerBzKbRnZflQYmibKF97Goret6
Y/KN9sUCxtQ7uWwqYatfYB19cvwXeRav7vJYW9XWIktJtBGiZNh3hp00/T3Kc+c7d2Q/e7d3y00F
K5Y0grqsnYow0A28UBq1z0npp/4BI25x/50zt0twQ925eWhz6xV6pEQGsXyjxvPJoeBPCvKqTkkD
JA9OxlPgcUIeucc7bdgaumO2hmZIUaP9T3SWgRosTv7JQa1iWv3r66GkSfahjnntxlBUPbXi+6ao
xLv949xJM2HU1rJ/lh92QMVfjgtBejcKY7wGWZBIwHO4jLeXs0g89BNaXWeJ5l4LjyqkYWlkkzRg
dFeiS9aCUaIVmgHpAK9EX1+75n3x9z029Otptiqu7qYEXbD2xiGhM+74pqYpGREQzDnmq+ium+zr
Ktx7+9q2VyEm8FX3UYJzQ7sDPJpW00RebMecvNqFffkv5JxCfyo5au0kiObe3SSfzClfDKkzH5sT
Z2l468xIQjBV0GMWi1iIIuYwDmueVz3hGzba/QCY+T0aUCQs2UN3MbfUF6wov+hf79casS30sMVX
pLrp9WByjkL91cwRjLZHN14oXKGT2I9KVgkm6yZxpAwLbQEN7FcMve5EAhGtbC7a9DT4pibOyK+C
LUD/hD2Zi7OzUWBGpIrZEIvMc2NQWyg2Po/O7JpMITGHIoEQdlSPrHhqsAu348X+oCvs8QDr7iV9
bKn2qczHdUqcZjrC5K0itm34oS+4iPMa7aY8Lot0rwclJDGS0e6blP1LcwlXyMWHYvy76rJtp5uo
+GrCqBZrzEBbMVQD/GSk7CWYghzj6kq5USVV88EMLVpnlgpAVpCMAyvvACmmUaJepVXel/gXWwjz
zfd5LYLAhea7bSE67B+lO6Wf+UBK1/2Km0n4mKpeRHnHSVgRkMTKd5ZiWMLQS7Ok7AxcX1cwDy8j
qos6XInVOKVaAiod/0WIwnV+8v+i0iAo5q+1dZYQ+qwh956syIzPVPKcUH2CcCZPd/LLd3VPDKNF
VZrMTP276gIhmUzuv+F3w7TZvX4HA4zU+4NNLrktfHVRe/xrz14pRMIXYKxMfFvZle2fRxceawgv
HNw3D08oD+BFJfAp9eYozTxc56M7/m82rHOIv+wQlEtNTqiEz+JLQ0NbYUyI+VC9iY7Hl6u1DI1F
ZX09F1gcMLSzSM2UbRPMd44U5xINfAXcKCNfYZFJITeB80c5PnBbqn2V0pCx4wgFvCYsykUSoKyd
ZeTxMbyGRPanscXM0G/UnsNMiXNyQ/twMe7wdXoG+qKFjH/SQ//q8qdgdqJlP8115EbOgGrd5Lfv
A7VSEGmT2zQzXLRRyViP3ij+x8JUgh57joS9wxpfqG5LttCPu8Vm9WEogOvz6bjuj4DvtEdSSouD
sB1mnU01WtVdIeLwF8gLiiaH47kaCs6/28IAZMFMl5mX/Fg1pkJdNldS0A08cl6lscXWqUZBnsDs
6h75PDRPdCu1kvAFoWrsSVxArWuH78iPf+RiISkQXj0LB8RfSffDEj1A2fSm7feQubsB/Zqw6Pu1
YBevtv7HbRJuxktB4t8twmOTL/Fzq6UdCoQwyIXlLlyuuO+aBLbxdEN+liqtJNvkR1EcxNR6e7N6
smA3yXjY/zSVKcBVRyuJzeUuuYjUjPAD/jNZ7VjX+1DSECc1zc1j6KXSW8nmBwOOn4Yf+SZIXlgU
U7+Ix7nGlidYBDA4YcOzE65oIsZS9hU1dPy4oehv1FXorQMSimGHABLhUTffM41a1brwn5zKXT5z
CDq1AY3L0RG9VVsuLmov7jkHhF1e9apI0XetEl/nDTysw6CSsahxCMgADhWEW20kM3uFMRGt8K2T
jI+m7/IVLMHwGgKqkoLcQatxJ8V8/QmwO10QADNLX/2YWMbEAw/aRd06WeqtRf/jcCiZGm68aTuB
nP2i/y8bxrwROJJWOZR4xfwi/uaQU/gw43e/Zhs6iTWGh4suahQSm+/u7bcGXMsAVtr69b3NJ9dR
/3H9FFBo0Jv7EZSi0oXyhXWzT3UTMzvAyYNkxOKG7vgl1T2wn17xs9cGmeLMhL6QArOD6VSyk0DM
V46TG9YGqUcJcS8/jE26bWv/1DDzhDN6kXJ102CEKK5Ng9TlxKmjhtWcSNMR8gRpraDJPTq9VITG
BmwqOthdiRTIl1fzkwkRkvYsfOnzrCiAbjSqzKAX8wiyy1stfbcOJstcNpESDh6kno+r5ai/RmrC
Cf3PDpB0mpO6bE2DF+wyK7U1+hvgTwLw0mGWUE5AgSFUWDbPVO6K06JNN2L31Y03BJZLFGXqFskr
JwSVlGs8T0092NIYwP46JurVWGS7940Vn3+YgK8CmYzVn1//4Gxz3I7ZhylO2/5B6LLz23ZCokVn
7SbMH+OVddJqnaE0n8vys6eKJ/o2XGJlHkPiitFiwooCZp2PxwrQSPhXkmHjYPekZfWL6qLPwO1X
O1RHvYeuSd4h8fg7PmxhN4Sf8+j6UvWj50GrZ2edHd7Z60shT+Rqv7CxPPHROezjoUSnKDqwptlL
JxsJRk4d+O5jh1OjKkLoQTiLFdFVlClSI3sNUdD2dilLKurvMwxelF+IadEiKYn8vvTfyQ4txGH4
Z1iROFRKrNa4sE7FTsm0mMCSdkWikZGk3FAXD4UHL+Uv4bbm51VKSdDyqaKxFExtaahGt73XC8Fr
xDDF6pXUHxr7DHznYF04oQ4GaGwUWzJq+3UKjv/aygwYvrcOotcHPDOG3G+tDWJ0h64mk40Jd3f3
xScFU9ggQtzkEU79tbqEdpp/xFnOGsBOA1xk5aUbEuHi7teZWnIqvs3MLQIIAnmDl6opWTSGyLl1
omYNhoFAXlPaTaT1GTiYeRKyc6ZQiVszZMYx0WqcHFsIO1ZodAcC5JNU5ILenjcSGHhEa/KsczLb
PrefnU7b3mFZumLh2ihWAxFSWowTOsN/6tvybc5+IqjLETzrw+4CjjkOvv0Tlsx8lH/8pXnhmsM7
qzBlAQ5An2wFvjluHEXMeRCPV7IyH/O+ddXrLToMB5U4pe+NeAWjKbawb4hEPnB1xAipP/wPKNMc
hWlbqbQ1ZjXACeE4M+mCtRFxrq2VWSTPxskAH1zRN5e4CIgG9UijAhEiqQWLpSidfB/FILJe8scT
ffCzbY+YptLgd7MGJN46c9jGaQpHVsc7Q7AUUrYs9/qF1jgmeKrBjgWQfXVat0AKPIYDCop/MKXA
JRQ2zoOku9V+oh5lJfs0NQLu/lHGim0IX/howzP5golkHrnB1jFuRGBoB2AMKSPS+LpezkW63YK5
csLrBD80++rULrO3wb5discE7gGp6DxhP6/iNW4YxRt5yUodIEEobf51+/AhDVZwdf55l/5wj7Yg
LHmtrWxZ5+dPjTWz4oE1DMAqjl/apOjE+5DFtRoZGPi3ZsGbiXm7/G6Ox/9DZ7X1sAS+UVcYk04S
HKKswuVOasDKMxguKncrdoZxaoKv2SD2ELbGQPemN1/rRAMcjj9SVFNtyky1JFYTIgbsXnZu68tv
2DU5w3U0NE+9DApmltkXDCbzr7UTefBa5KtNDJzNPhmSB4ljhBU8cmhRds2tjPOcagAUs5WnI5Xq
OrkDbSzVxykiNF5J0LG6u7rhupwjvFjHTiNOrsFOERY5ES55s4zF4KohhENZtOKcfrTDM4xkOGu+
f0kOfaNcQ3ujPBuiiU4PuPGGE374VaOUAV9WYH+SDmSvqQ+m1Jcv0EuVCtJobBkeA4+ekzCIr0fm
4B+Xx5yiMxvUaiwlfKPxaFQJRSLVtA5pg9IcNISrZV9/m3oQJBZY3gDQPq7tQf3ka+CHiGyxgyJG
+GoVJUrhxLrTBSbaGP93EuGOknX5/B8NDjF/EM4PXp8n9qIDo/lqI7Sv8eyrvfABMKvfyItD5Rpx
Lq+utuCYZACSvo8sl9a17OoxvH+pIy/ihm9lFi4PcsGQLMJRLihq4RNKIVdYhDsDZzYkME06zd4D
DKgGH6R0ipFTLrrSxkOc/M70yGXD0ENOfMUc+801FBY6iiXh2TIFIu+6qV75XqqvFsujMUv7Gs4L
WG9uzM20Wqcef/W+NqQ/U695coPDKOvaajE30wQcVAERAyAnq7Ai7czDOHOm5RnGNGQtoBdXlMBG
AhI4tVxX1ibHUVpHndWy6k2Dqqz03Y2eTYOYLKgocomh8Dwn/YRCjGeuUE5CUJ3EET0BBR6aQ7gH
+wm0TIbxT5+Brvsj58Boj6nFMABgXWVitr6Yvj+cTRbApQOx/L8ayFcEvHdSVX4vyGP7/w+KUB0E
BiQODWkFhnWr+DBqUud1TFfcN5+m9j9BJk3b3PnyjMbhSuH4m6ByxwRfuCksB+sC3WYU0DxB4Ke6
ZfXfIvjIGyP8awfbPCBHUnVBHMl15npBrq4GR/KMkDi08pG6Chi8j/5WIOG2k7vxCAvuNidDSZqr
UIOA3Jv2K7ooqR4dRvb/dx+m/4NrNIhBYMIoGkynLZ1r4skOQzd0QIpovfWFHMF8QwARydy5wYLK
V1yllBGPbW9F+gCeweNjnLh4p3MgpQdXnnJSuv0YJPu9lztazP7TYSTKlVpUPfTO/td4H2PBSLYT
wpQy3VZGWnB6Ifc0NKyi9AF3pbHTrIJQYHFzHmQppqVz9Go8VjAqhWQPDpv/vvnk6iOTPsnhzWaF
YtR27zddraqnB0oBRagm8jGKBQWmoTMCgvWpts0U9FHAWVLNS/l2j94kczpfQ4rYz9ncXWISD9yw
vR91rpRZKX3UDFys6qL1iVDEOg27h4L4CFvdvmFUg7cI4SfqlA0JLTv55qoeYe8MNmqj7l9sZLxm
PN1agQZAunMqeV5fGzLfNHnmO1hg3wM6PA0oq1QawjrdvgYeIIwb4vLfHHIrwdP39qeGdVzqZhEm
8PS4CQFu87ZclTHl8Ou1c+FLEZXrYAT87DwM3Mn/vqGhkpxeXQ9R371O4Iqa4E31ynx2xIaT6FJI
dqIUPcFWSZ/y7ML/l9J1nsO48742a+8M/1eNPSkl6G1MevcKKxLPf+CR2WRojUodEOpyizvekNqz
Xc9dTZDgNheZ90wKE9gkmaA80z5UPfEaBFCd/8NsiEe9D2pW3TuHNrBo57Tlaq4CweLZZQH+rYLB
KDF2ETAuj4tP+JGjc2Tz5HhixJM8yK9U1UOffBE1FrAeooprpXhxtOI18oBJj0HZp5CkKbKc8zCP
VJE85V8P2HIWs4Nr5b3csKtlQ/+13Zkgs1eG4xctAMkYP0Yt58g6rapAlAPcgof37nZKomUXI1Gx
i6cl+npCKufu3Wa9uYwXZlrnDCFI+OlZiqH0oYzWSjart/TD/jyQ8v1VQdu2JmxXXgz1vNz3nyCm
G3bW3jGZ758EMKFjVcurcF9e12ll7O6WfAvORKKodzMHpL6yLTZHj3/D1c8LyWHIX4L6G7jjD8d5
6ZSlNeUTpsgcOQEHmfeKl66rW79bHe1emX1kT4BcETJIHLyxlR/9ySExGJSrMPMGWMhOYobfLLUJ
trmJXsk/eULK/aKko79n9RM0OB7irWV7F7WG28yISTCO711W0IXY6L5+G/9UTdl/PDkmw6B4maOq
3UOxKAGKAu1jSqxZmgk4OBRkYFEkJ/hPDNy7B9st5D8GNFkexfT1KqRlwuKz1+H63AsJKsXVGju3
Sqwb8cGNUZaixeNTATNFLq5J6DiyQXvxsBSzgiSYq4mgGc1xNchwVG9IwlGkfpufcR5eZNTw14Sw
yyWIWA4WHbCeZecVHKo9rMDfzbr3r6JH1Gim3RIuf+IM2GQqGb8ii1YkWZCJRlgBcLTFauUlfUwY
v4e2iKE6gEdSePGShZy+wsAWuH7EcIXBGMrgvQ2J8Q/Z9jVvsvPgU9nJH3Pux0ZYS4kGE0ERu7zk
vw6zHI5O1JgFZeK1QnIW3hErAgLn10VeGXOcPtgcy4yGtSOXkLfOtF/9BOR8JT1tTmvqK2gcwHbL
35eXfRQibdZQgIh4f5xcZL4hD1KNztO8Dhrj2J0LDp9u09evxliTD4dusZLiU2FL0cTVBfGJC3f2
o9VmfBG5J5IqFiNtj6JOcLWPXfckodhGW8oeuYsVgxqsioWonboQbON5zy6i8+iYThajeZ2QbaFO
frd+bEZQfaTDVPKsDd9OCaqyD5/e5I+eltZpLYg/AcgH1cFXbi932r6mF7dXAVRYukXgld3f1FAO
eGJi3fkly3A8SnYcWckPB+qf/aCkcsqTZuWBX7UlccSHnt5UcKYzVfBhvlpTX9gZJO6QjIf/7O5e
uMdPnZrcIzjpC6ChhoRj5Njo3ZB5SJpUxsUVBBOtd5BAhpylKoszQf4ab01XlTSalGSnBYA5rUKw
nY/Yzl1za6FBzmHRC1XxKTLu5gLG8F54mJAl1IopXtByDzKb55xAwFTHcQrFTJFIWxyqTpJKMczB
XKC4U3efFAbws+1jOonKhtvAMCW7WZyriF5EkZGhk1E/Sz1ugqEB+n3wiPKJvPtT3xnS2oUWALWC
HWJiQBw4MmCrD7A1QD3p8o+cUts6OymC3rlfoto+ikhDoBJaiZYYnBQpKhZquFEV2hvtL8nB8X8u
uL0K9q9u2OGj+S4KrjiIDmVGdX05wqS+FMN8TPzzG1cFakK/Zzh4kmhuDERpme/r/1EYMP4LxDaj
EQRBDPBib50n6wbxHjOaxlGthf3GxgNnqMrvrVfpnz6Ni41TfPXMnpu+3KWGfNxUlwKpuZzvQvye
dXb5wTXzWHVmDOSeE6cPAYScAD5eEKjtNzR4M1LgKJ+AMSsC6Kv6pOQIVJJyq0WNXFYJV0bV62xA
677gcFciTgoABMQtT4t0kBB5ceVyoUBrVlM860PvPHBXdQlV0rcwS8ns6SrFctaCx0F5CEt1J6Lf
lqUypvB+fkS4yOystRQbyUoT5sKKuRlijz4AGHobw2yxyOCmX2n9hxcM4qXGg2gEfohbymQz7HNH
hN2jp6XXUB7pNO43Vt847PYBxHzTuGvUy2qyjUNJas1uOGRun/kVmKHiUDjtyomE5cYb6r0sL+VF
zXq4glaxS4ZDOQQBAC0Q/SLEopIi1QjDfinBxDonsIXKQaskWiZH1ZyCzx4cqgZSAsDekzNHGgaj
zl3OOJORGYZojHlYsqhIlefRht0Zz6LGH/Y+xF/CSprNX5xbrn3kY21EtFBduWZjFSf249PWaYPp
lQMzuKVbLEQYBsbeNjvp+N+t6qQVhXMDvFsoiBsEGebJjY1Sb5RrChf/8sEv6eEAiivh2ib9O425
dzjcrBIbhAM3N1dRJPQ4iHtLeeyCmgKRyhjntMpY9fE4rS2XpwhEDk16vjyDfioSeNgB+1mgSel+
mzk2M+nnMoKcxTOOCLcY7dqy0wdtcL2H1szgoloP63wiDqYAiQsliOivSPgBGJrvaiYErLaqxY0Q
KM8JdGE+3gxJIALoXCnRoQ0vkLZVowT6ZiugH/pjpuRuaLz1/SFBMjNBhHqnk7oN+tKrkcwe7y7P
rRwH+fckBqhh+07sjst0N8wS1rFVNh6mF209X0u+0Y4SiowLH0W5IWI2jXe77o4CosibnZ7aSEJj
IitOfyURLzsQB2wNXATdt6Wox4lgP6dXAWVy7NwvP30BDL+t9iD6SrtEkTF2m+Hi21pm6hpBrXdu
TmpHWC+UXS1bioVsvKi+46kA4wg3VYVIP1nlOiyGqqJKH8lCQPd+JIcGc/ePi4yA40BA/uvZsYmc
VlnZ+7U4/YMbc5yhYQZzIPGNx/A1nRMQMiHLVUsNPmMwmsZhobzWneiO2DoGdqsxwjsCfAPvNJJ5
3LAH+nl5QMWJsqvuDNBJUyU5pV/tcFdXlh1dHebwNmjA70LkDEPHKd9eFdEYkPpNTLhvCcBADzs9
8A3nV4jr2I7rwXirsc8GuImlh9UdjHQ8sDqhZoZo28cUiTKatbEMvH2DG3d5STJsgsKIPNFDimOA
TzEyaEg1/V1RKjuVRXOBWIoySqsC0pYFIDhkvPBsS9XUKV03pyc+pwsm18pB3FzYWT0EnoTPZUcC
rN954J4HoUSgfB/UgGldSlkdRiUSBc08Yjo7SsQaIn/TfosoUAcnsS2NjBXVZxtL0FDwDKixwVzQ
2DnOalXRUOmVEUXWtmO1owhL1woCSIBbkgWLEnyfcJ+z6WCyh+pQM+SlrYv5UEjoVfIAl5N67Doj
4Anz8U4P/BNjkv9uB0/f8nGyvyfPgr3y+GhfSkD7LPON7M9nCwzVEgF7NHNsOenlujybcKzt5E9n
eE+0/8bPSKADQzKMR5+1uE8eKB2vBoi2AFXlm/ViVpkvN0uIrsWXYCDy2Kj5NBCBbpSOUrR0CJiu
J/pl+Nns1oEYKFrZKTzm51H3KkVEWc9PaZp74iuM9G7/mwQRx6KVcZj74WQqVFXwX98U0eSrrQd9
8ZGFPAFcpIIpOXzFxPVf7B9Q86aR+UKAyQewdcwdPgRO1RcNTdlxRmLoJZyiPPuY4k00WcPeKZyl
5bq1lhwzQyBUPnk1acoZsXhYc6E9vq+MbNxhTg/VEVOIXTSSRCIZN2qRQBSsr3d7qgAV+VNeRPIF
ZhhxIOxIHXM9MZKouEnsLYrJOgp4AFsIxfwjx6hAsQ3aC0rzfOKMxOAXq1izK+Iqp2pNAOSw22fF
M67mvclKOL+lun0fpIxTomyF1OKIDRYEogV9Ib5hLE4eLZwRbUIRWVRDb99t2T+oOtcc9jqUrYUC
DJQUNSrR4glxj6FYLk8NvMXlLqxWY+jH4WldOY+dLINUnvI0FYqqwpCYdvmzGE+X9aOxXsJ5IIsV
Kd2HnASzwtSML5kM2+6VDMkGk18YM3aZ/Qz8zZBIcgudtxB7Etu3AyrVZWVWVHZ2V3sAuF+pJsKZ
y1BWPsFsz3BTCE67NSz5S8u8IBr16b99/1b7SqqxVrWn5ZFtwPaqDdSzuRYaMhe55PMmReoo3/3t
lup8Kd8SMHYJGkulTRKmwTaB1x2UbXOtrAFEkEkXRpYKBpAx8ogqAGWLc1I/OTr+IqzaneRQaz46
hrG5LiFp0RzBA12Jx2aWMxh+Es2+l0N5FO0wchrQJTpD3J2hcxgx4xDLK4olklBp8ZsZdshavVBS
cWY/Sc5lrfqzY3GESBG2MWXANm6xB+kOVInVwxZ5VOf07NYS+rnptT0/6qvnhVoH5Wc5wBeVsw9k
Z4/zDM1mqZ2sIrsdxaiZMb19edbO/gsVksxVir47F6bRE5wMQmKnZVMfJVviNFxE4QXp4UFWZcHk
N8emdyZ1WdXSJp/N7w3B+zhRJ3XOEAQk9BlcABwpvsSlXRYw9icnhOJC4sqmdWyYOcFnw0DS24p5
NMzKAU9TIehjl3Gzuy7+LCJsLD2GVnEaQAzVKaWGw+kfZNN7gosEpCbTcRwMhHTqXuerBFoKGd9A
7uoJAp+nKnPSKFkZMFIw8BoGPU3kU8g7Ykb1wUHTQqei2uSsbI0po+pw1JaBzanyniJAVERJYtDe
66adbi36XUWg20vC9H+r0uhw3S8xfGEKpRJ9ey4MSIg+9ydX2csl87aVORtuZevKH9ziYUnElfkv
9aFUV6dlt15l5fgXkc/hQoauuxixWEWeJOUJf1RSaMTNdFrY9lGmzEzW6LLWzVv/XlK0Cu8g176s
zcd9EMr/wQk7+4GuylHDzmafZJIoPIB9T4uAR3oR9P2UGVCtfVOCfLoCcKXIdEp0Wt2ONDBwsuWT
oLSqLJf8LVwacen/5SQFKsjolbRHICXer2gR0aEeNTxDEVWn4Wx7EXiK+F8UIZ5WYQIfJfToI8XO
8Q2uCeWwut3SZFhHtX/GJ3oh7YbOHJPrRNoaKbLSPQjMkUt1FFCjLQ9j6yIA9ptii1Qwx8wijU7D
5kWJ0vLOtBMpH+GEUE60BXe1r/sSS3LGuwApOfgbjl46vwGPRJfkUoyg5ko6qLUzKPDQkTZEAYFR
5G6SFqIsMthlytliRa+LDpkSRNyi3o32zA2IBgxrVWiA4zJtGp9FWnlfHELcQqAjuEazZ/nXI3Mf
bkM0NUjoea+IuDCU1ZiQ45r15WVSBy10k+cYat6Y+Yosutxh5SP6IpLRPF+fg1ixz4/580U+O/f8
GjrelaWgRgnzF1evEph9iOT08Os7dsCzLU5FHPjIz0glZHjIhV3O5Hir+ICu7XVpLsFzwHstNRjr
ir7LW+5vApDTg5NL2OJodzD+SRt9tF66k3k4c6KL3ppoiViPSlSUSBmveD/NTlob+Ai4YlhnAhQ+
tc0qJRQ1U5CO+tS51EPIZBwXipu6e5RYx0XKK/N7fOrOnP6BSKmb04j3z3QxsHoCacqRtIkOnovh
t/9CMjRXYk29abK2lwcQW6BU1mzIw8fwyIedLXLQVQB65YuZBhRl+Fnvbj3P2lRIex1mUgtLGcac
OvawESLvTwnoh4nIIaczaaJi2jY8fwqOy3kOfQ5s7ZlPHiq64EkT2TYMwiwoOOFOk/goHnZ+/8XP
xU6ByBrLthkWO9rYLlUeC26BTzUmAjSUsITd8woxxEz67mmJzN3hAU231L4rKqtZtLLAExGHDeOV
0x5wP2RJFy8eTYme/6C6FY3j3a3uvpJTmCBvnqn21HI6qRwGihOcCQMmGTEDZOkbmPNZ2uVQ+yyf
nPR0IgVexQgpcTPfvCY3SO3oUibfAvu68ZHufd9w7hgvo3PSGWcQCqVw6Q+OJSOb15Q+8AEvqD8a
mQQ/0AcNwgp3Bq7nwCt61Ln2vI8rbCYEm+2oOlvvmIygFr2593RQ5oqb7CjZm+SPoAnF5evJATJd
TSdLhSvck2UHqPpXnAWWSovDTQnKHsevCE5+K3tUB14uRQCdZFaK/XA/Qo3xc+DVY94de9Z212Dn
wLSgdCInzSDyVw0j1ZZTq8L95C+ZFQPCOay5VaMKvH48flzDO+ZRR5QWM+WLdCiVhPcnhT6ldnqu
REIskJj5bIA+kEC2ykiG24XcsA4becrmRhIXDSF8TI3rOpXPQOvmblbtDVOnE+x1Cufq3rrMFZgX
qNXf2xdUH+iUoqIgr/QtETgRIMnVFTzU94W42Vuma/BhAedmaG2XLsNoYLOkqKZu7Z63ghM+wP4I
uX8O5s+B71TfJhZYL9GjDRz1DNRNUGvUOmGRr9KUMrY279khV6KFzlzZx5EtkpanBUp8b8eCL1/d
btNytr6q3LIwmh3PKVR+ecIqpca8bHb5fmVMA7iuOHLw7pplsxuKCrFlalZlhgm/hB56QYO1EP3c
T8Bmr2IUmNg3cF10OSLFMm+oxfoY+Xr1NUEUxiLPs9iNWj3TeQ4pVzMGcMtwQdRkYGhY26ABiaBk
yr6G37inHo2FcNw01Xixki6WBnkprwxhSSSYpQFeIW/YyNozVYpohA90wBaExJ8PmSQO/aD69HwL
ptKGH9VPqfe9J10LRyWhK3Zk4avHRevrXjtpO7+Ri8BLhOOZNha9MNF52AyK7e2to409wbW0wiY6
kGmWsCssZTZJhKsHoM/6FFFiZpBpeINpkIT12MpE9HwuMfqA4L8CWIjefHAPZk0e4u8yRgCXxbV/
g1XN85ITkG2B1PP9SpiAN2fNPAssbCFB8vO+umtLz/Y1boyNIKTzN6OU3vlTZP9B4oc7RU4J9S6P
Y+t8UpRRN5FCC5MQu5s2SctzuLolcUOjW88M61MKMcgG73EX1/xoW3OUssil9C32nlqSPZseKmk1
5ryR4kWrGl6VFFkej/DVMnjvOnt20GyzHAV6SYSKIv8JmNs7HhPeKbqKL0/ImNCcmwRU+49LIP+d
9U/aAKGGZZTpAaqwrIbJUAoKSB3JKwMVxuBExsanzGZ1XJqOKOwuGfrZWQuTm5mdvNsZhxlBqMLo
fI2bk4uy3yaBOgkhr3AihPWjubWV3jR6TnXOVj6PQ38LCvDw0f1ZMPPi+0nHb6dlSaxwX4yw01yx
Ru4kRBvK8nnJ1tJ6vnHRUu3xus2GyEouwmyQ1cJsZIYtJA4Tnc41Bgh6/Zo+G4NJ92rRr7pAjVFb
HdJ08a5YUK2oUuGe+rw/HFdgF99CqCW6gH9ZxZlRwGcxbZwTxXPfKlEdWUQ7MFKFvzm8LE6SO+sj
BL1b7FbhsXuRq86278Ld0oC6iZgNjGS1AK/mpc1hyvBP3k8DWIqjZ//4ALT6RTVy4WOgeb3U39bx
CF8EpPSsiL9ArDDq2k0K2Ylv/5OV88xA+R9zgg7tiiVXpkdLSER/eziZdWSWJq8gYjWsvRI0mlL8
EtclYiBUCKCmZ+kBp8BJVM8wZEUBa+59jyXoQAByFRBmgY8F18XXgwV3pxITlbT6lg0LXJOh7102
gU3HMWfEXes3k3WSYFzeJChKBEjLPwfgBkLl6eaPlbc8l2qWupPMkMsLaQI7c0Gevt7UX6y/3YUy
PyfVaKGzw/hzU2jA55rWmBYLnE9DyK313CB2dpyXxdsXhuvnX0v7TEozrnUsaD4bvy8HiXYyxIem
YY3gnyAq9CGqntF/1er+YS+UokH5MTOL8t9wC0PG5PcZCi+T5U8y4xz/BBqlLNzOH5C7HkI1BP5A
oBYT0bjDBIdyIuOARgbwnGaqAIPpbTmLhyTBwynwH2DaJUXb4hgfNNBsknSMNdJO4FOwkOMNbnvS
1o6QGrmVRdP8R4RvF5QkvS/IATzsOaLMUL8m8RV6PjoB5zhg0Ahebjd7C8E0prrmTe+ECLUkDxgA
TxSeohd8lKwvmGkv3OSDSb/X7sVzsP6g6426Ei7WAvFjE8Aa+E971qrhe6tTW5fv6noWoeMAZyyJ
pRnT9CGZFuguv0UFld6xGarsPaDgBYkowtFkgpvFhGXpxTGxBeqlVm3AheV8R584jdAG6fXca3Tr
0yHLiy2jD2M4Auu9U/2JMScgy6dAPD5NlIiPGEelo3XLY2un7RT/meGhEZxs+qlQR39tRXumztNF
Kwpp+wy27NuBYxlijzkTs2lmoLGgf8lK2McqMoVYuDWsOwgNk2UgQ/4Hg/uKcbs4ULO31QeURhi6
5l4WcPSjFXMG5sb/viSpXyoLGai1VWOlOoxXN8ZY7c4bTkOIvlE8lrxDpePs/I18zG+t+/go3YJ6
BLLmN8n+lcycBOQztuxgbFUSgNq5bLbSUilczcLwQjYUEJT5NLowSNjqLmKRoT3Y6kGKbO6BkakW
PWy8E6ruJWlwPJx9s9iXA78NcvlSQXCM/ptn43hPIkMmcNxT14f/0IDvesZDl9OttFbYJ4PVmgVu
AwikMil1fMN7/p/qztk+F+tWvzKB1qnLrTZx25dh+Gk33Wj5gOGjZvi+nAy6pHU4tYpxMXI9BcH3
/QFZTJ72SR12lRKsG+PerhFXq/xxn5wUcqTbu4VmLpRRLPsqfb1Bqi/M/rHlrPdFPrbK+xYizJEN
i1qtk7c7/yYxgLU2mWRpUk+5M2SPbMmhSvXECGwfStae911NnALb4E0VR5AvO8BvrK8WzPkJibw8
Tf22u4lyQwWbVh2KQfNof8WK486qrMoCxYkuCovE2tJJ6Ios+2eUu7xewH5rde9WtWPZKS+FEGjD
do2zVAikWhvRBuvHjgaDG8mU2CzuFGkcOgZ5u5j7RUYs8KsbOIqdy6RS/R6oLfmtmoUMnjmFHhoz
hRzlOPWlv2m+z7tYXQlflVDy/6hFuRSXwuIMi3/M2Q70F8JrtBWkLjcSXlLlmJEcWIsdEzCTFlnL
d23pfVLMup3yAILCon9v9dh7SpQUCiFKEdlCBiEfXqJX3bOmjXOOuWAoTyRxm+kRFxTstNsmUNkE
pQ/hTojmQlj/ybEkuwHtWUQuZ+xUYlaMCFqfOSSf55rAJv9v2G+a1WzVJ7Hx8LqRei5JfW+zM/wr
1RUozaR4c06OpgpoZM767xy9XWVAq5iwoavHgSIYmNLd9BLI9ZdB44wjO4b9fBfhuthXMaHDktCG
Lz0vl7OAC3qABkp0KpA2e7fGgPwiMcZUYYdeVRVE/nhxkve1LAxi9PRyGxVAvgnRio6SQj/1QqhE
5EJYpsmFtQyjYGuBsJmHKGBFLL0ZsthIxVCviwSGNX5XA0KgPZEUPquOptNKqm5rA9J4pRst3kZ9
zRpobiAHPzTrNwNYyMfWN4drMopWZbNoVnbASIJPOSvjI/BAMnOlWRQoNK2ujOdR2y582+GVUnlT
6FrNb5u7o+nLh+nWkj4iGixqlyymsaU1diGysxFvfCJrMEDPjzhCx2mbnSSzPWWtu2kF8k5C2F08
Ee2EEdJCj9SlDUgn7Cfa78IXT+8Ww5zsPZJXOAWsLUXwUClkGaSWIRtOFXU4l4VSNS1N6wlruYJK
1QxW9wUrp5HfFhqx1bvs/JGrRwJkBH3kUn04r484/kQvpeb9zVWlGucqJAjLeG4nJGp4EkXFsMTS
yfgKprHWRfL+hXyZhbiY/akpO/hHhRCCkLzswxocVN0hNq+0d3BCA8adJorS2LaSHJ9Wkdhe1vKI
uAA0kQypkAkaDlHVGHE+O1aaJg8A6sVw24f8Wx6YS4aWwzeIFl+AdGCUr7KTFJlkmbdiD+dVZFuc
gzqA0pksviMJaG53tDeusEfOtp248GO9eIqrV/3p/NyRqrK8Sw8Of/8PRElozaPNSEulASuMO+N8
j96FYVf6g3Z6gYGHHCdntlvOkYSea7MkViyi1YoqDZHJz2PieddOYq5EkQwzdYn6Z3p45dkxIwyK
YsQKzLtPiTqTltHT3q1A0ytSjbW1BN5GdwHzXl9Uq30/2M9yic4hI1vt85E17qtbDDZ+I5HHa17m
WZWYZmoNV1P5JoGmA3XtSgB/TnHcMOo8KCbwq1aMZyZfXk+xn6mwjX2TKx8fnmw+AbfMi9YRI3SL
67dxHJV8s/53yBDjRCbMfc4RGDSb7RPIT1+7STnE2EMs2N+g1GU0/0RPgdPaMH4ZPYonyhszTt8D
rvFRTQJt3gHsFwHGimzME5vwG8Pvem4vHRoDRYypBBuRL9VBz+ZAwZTJgf8nfHODXQeY4XssGKJ9
mIjV8TXKcGj3kNh+WuZkyz5PXP8dQdV3ZBXgaGQ9lsruzCwK/mn47IHI31VlrUSCenK8akTll+AI
wMAyV7st+QqSragEpNqMFzttz7NH9FK1o8kY2896AoB+BRKa1Ib7t+HrnwZsER1g73rHo7f5tA6D
gmpCWCEZOQ0ZpduF8dhVGsGPwxf6cUA6wmXeZD7O9aut/qT6kaydwgC6y4kHqQ43TfKsm+CSiXmJ
AP5u6jiVJV42TDo2VEseOocToqilSbwxZEYsJT3c2n/IojYu38V6q1JSoJ9wv6/TbWzw7scmO4Ss
sBvX3jJozT8dV9OXhpheky7tytnyZHC7NVduMHhnd5VucqaXkMg4D6BB+HP+Nj5oLJzlo6NGkvnU
ATc4mb+Uupe4V0HXVEN/pj2lT28FyJjNnDf7hv6CR/pwkwBTnN84rnuzXkMPMBZrhorfHwRCuk+8
t/1iHSUL/gmJwORd47HKpYO3hElCqb8UiRZs9lqZ38Gab36r/+qQnfbiLgX+WIEKEAJxbgMgGCDz
pTpYm895gryHo7nrHb8vKYrVP4EG9zjeHdQ1Npskda5Yqjb1VsOwIkUlwRG4VaEoBGCrBB0eBDyB
SUSIB1ZmGXDBBepFPPY8Zf3y+uQbNWmEoRtBK93PAvEpUaq+4csx4PRReDgtPIAKv3Qmq9P86kL3
v8SNoqUvKkwaZ/fgBBDAjl9d51bwizCBKDVfqIn7aHUiBVmIf03zDSa2vPnUdU6vEgcdyKved9tc
WgC60dWldQt2A9ZhwltoQCLozPI2+V201x4pQM8JpzEfgRmXO2iOH7QUvswaP2/0yl80Wy0s98hZ
gJC3jjwa/Blws3jmtYK3ChAL0YbWzB3RIRhKOr4x1YNkefD3jc2DcSUrOPGblLlTsJIXkwttYJCR
fnxhJalnqLZ4RRGG5mEZGFXOm72xDaC4ewrxyWH3R/MQytCjcAAvHJq5faoAzvpD4xPMt1VDmqXs
JtnApUjKkyva5MsWqQHP06yzCSR3/4L0QsulnyFOm31LKV+9Fm6cjog21eonomI0zk58Q2iNuobA
P6MrtXoHD1zPk5qUx3RJ682agZAfJU6E8r0cl8ftwgPZj9Rk1mKkIVAFdAXxHFLzPKyCvv71Wd7o
cvpawbML9W8gET+SAj73Youd7Jgn/XqP3YeSTU5+6mkm8rUmpZhXFRflyfnwpl4MCs8t8IYU/l4+
dtu/DTFb4P8nQC4hSMJDLAVcPn8sch7xn4HuN47pFrtu/zkG+5HO7vfNw95irk1ulmXpjvXu49cF
Tqvsn4H9mNDF7qLLAEEusI1PfGyHWJvVvAOscra/GatxPacUlWhUM6uxSS2hjprgUV4S3ftaLWA/
FEbStAoKdj88fEGMCMDWMOjQZH5IjaWblQzY5Q2RXlFQczfmqcvWQSwBSfauL98X4x34XUA+X4Z6
r1w5Eu0Go9SCM8KVHqsurSdymLO9CWsNMdJHF/eaav7JkbErBarwTegzsW2H954GDVogGph8HwP5
4tDRASMEP0B8d2rjR3bD2lJcD30vtTsfYcRWAKciSH5IEoZEWJBIR0dah6z9x8egsbVVP1qY47rD
wQvSpOObUB9uyc3+EFJBNh5dUIAiNwoOY19k1Tn1m/SEETpXYvR76Xk4ihyM1Ga741PvA4qMR/pg
REJ3BKXqGZ/5Lr4ecfUgRuYmdlblNonU+leAd5U562ViF4qBB7VBv/2bqbbsZAVqPgex3utPBFMA
3PkG7U1TJEvJyK0xPRtNan9MKRUQiaAZpwF4dSw9zGfIWv0ef7b+Apn8Jsp5uAq+mAuk4k3x6qj1
VeNQWxf00/jYvU9c2yws+IGVsUas/8dWWTcwzBzD5Cn2WgmO51bLcblvWzEOAxpJaHYwxsi6QSJb
97AKQs4ML2S3RmRS5jo5oKIy3R01uTmnUmNIhQyiYL/cJzo+nMlijnR4GLPBKxJAkL8pBeTPjNn9
AxGIVq8IGi2yVwkXuMUBbSm9qC6oG0vvL2sBtXcVTAyKehEITve0+LDLcwxqA3I98FGLGuAWflhi
6eUoPFXwCxLKNj3WZMYoUJH4MyE80QMxFCWzbXkZbcu2lPHJTq9zwUbp9z26MwaS1QskZDvwR+AF
Hs3DcZXOJDrH80FiKfx46OjPBLbyzOOOtLott0hnCguN7Y3uqJN2z9/ZfpHPBhovB98Tj2GMA2vx
NQKBq5uO8L7Uw/MOEJoBbpUPnyN/0e3LIl29aXtmv1RX8L+oaGoZ/91aHX3O8b5mRGjLm2k4CTZu
ti2TIFQVDXPHuRrp9TyYGkcGTmRyvvNEuQTBcNK4aT6rm0LW80bETAHhkRuhkRa3dhBS03lV+/dr
zhEwUDnJb4Uv77B+p9xdndedmT77yRpVgVNZP9oP64266hU23K0yx0wEUi3ToHqFCjE4kJfzEeVi
WThGcwEtOTDjzCl8d6zoll3Cs4p3vJVVS2UKDcL3ZQZlRpozXEDMcZRf36dYA8KFnLGBhQdLQY+q
SfMn8JAglZ+a1NrNk29t7vDDIAXcLCYP3JOPcXr5BhueWbpUTTHUW280/1ketydSotwaRR+ktUee
i2vv9zvNxsihmLjqW26vkjRpp7puJlHgKQq9nYhFZhjOrGo/sZ3LKxAiCc23BouvSbc839Ey06Vj
f/OU9014/6XjEnZw8DsY9L44KluUdTGsByqt/A/3ABnUATsm3eh84XwT0yXFJtuICj+0IEw+0q14
QXzZ7uipV8cKgQYcTMTgTP7cp+d4Zia908ndXKNPNcRh3temLTMIMLKwhd03oFQHnSEFR2NUbUWL
9anIQHtmqOZhyASKjxeBmSOCHDv5oGRcHESXh86pG80miKfmU8eiYm7IOQli6RSWtaHOSwY6zMMS
IjZdpogQ/xzkkFqnmLDZEfAFk+dzrui3hl8G/f82WWp5WpV8dafbbzkuS6lhxrALcVfAVSxPQiiM
0ELI5pHzTGfPsRZifuAGJJg75W4tXV/QDnZP0Vhonjf5MUlW/YuIO1XMsVEDeK3cx0cbJ9yVUucH
KQhNUdpZgyTtAkTzmh+UKpWTJ1Po3xWmiT60y2R3e/YDwFwgojRVHkm8ocbYpaENHUJ9PwMxo5pl
UjFr0+gKT5bJeUce8AcxDzypbdRx9GsSQkqKio1fbnUQYkS3vVDYGktEqkVzk1DkptmQHGSE427d
GuKu3GZ36Yi/Sz/GnG/KHStGhT/7j2WgVGo1CEQaERo9lHQrApmWWdVJiS/6s/3KCP+7LVtNG7UM
HggspIIsNPkV01TS5zdmRVjhnQiy8xCsjstSnBaVVBcPBh2eFdvC8/CX0aMG8om+uuGzgDSYfRPz
Gn+ndJi+iuWAw0+afjZvU9fEcHVMJ+ZZ4Kc8t7Ug+F172Pveg17YzmaCm2hKEcz4iehKRqsZVeT0
kA4oQ2H2cfh0lLR5frBtZ1d4bQd/EmN0OxQV7qIvSfrUyVuyRn2kQp7gMRv2P3mfV8RqESqINBzO
2OU6ZCebfO572Fl9qbePR2HQVtrsSwnYg5S3/OnxypOv9WN5gcbB16O54j6A7z7I5z/dDSViMRBU
dlTexHUA//BYKj2JlSifzd9u0jb7rhtsax+DE0P7bBV+eYElihv3O5JAq3akFK+PzPrfVmd0Tk26
tZMsKbYi2XKsb5NVEyyegNdcibQb4p/beUhaziAxMvafiHubxTGTtvVwPCWrDsazDPogTIQSYfTI
fsMSVxUhotUpzz9aVNdd/L9MHDNajsIIlC5fodOYF2J1xtAcmc3mZyWn5alu4nxkO6FUWPN1eyJE
EhfKOliUSQ8Hhv0O7Gw6/uUzvnDViLgHZHZzmDEo/21LPHXLJ3nOO9e72MWEd4V/49mz118LIBqy
uOwVVtlA6Ccyc89b3BaJoXMySaZKOTSv/583vJXgvq20f81R1iHpCUCrybYD+V6fBXdojZ1IxQCl
EdRQizIFr9uTgUqbUnDgMh3WaXYY/qIBfQs9bwLsmmMCjtGbRKcP0tZv7Kooc6UCHJ9auLz98JxH
7WdKNrgiRP0cLqdQUU5o9pS7f+LIFi0en8wIShfotEJNJnqdNLiDJRQLBM2zsbHkmAuW17XDib6o
m+jvTGb4H+/nL3tZKXvWpWmTFPhkgsoMha2rhlkXHp7C/VVS+t4AkGHLGOX4xpc1Q9/ADIydJrHO
oLxwAhMbQl1xVxv+yJ44GkPiUNPOyz4AOF0Xqi6S5bIPislGulFSaQ3F9cpFIpZAQOWdBITraZXh
m2BeIg4wD7RwMWI58Lt7XPL9DJn2jBqcj5blM7RJxCTpdKEN6/DmA237UBA3eVArZM/jZsCtmr7U
v1VfAY/aVLgwgrHhZpZPmNMLfbro7OPfzaI7R6ZIRIEzzuIZkfXvTGRWMc07z0js1tfGn2c/9AtX
ghhNvZAF1HSBVR6nc9dMjxO03IsmyCMJBNwXHH1l8U0cBDjQ/BSaJMOg0fwGR6eb1Q7piaiWiRRw
3OJyqY6qUcmM7nib1AGxS1o6xBpTaIwOqtcI4k1D4esRffv168c0ECCeYw83U9WFJGwxjSbt+boZ
2fCGnnBw/vPjtTwqHH3cqPpwbdUIs/stjeHGU8RMUgyoore9tMi1wxwcyFu++7WO/0mKEDMOhtqo
cqWp8lWZyiegQSm6hgGzUh6uJsQ4JXca2tcOICl2Y2ODx/CPOPpEli7tQ0H3+Rk62gZoGoCG7geC
HDglIleQp8uYEMMinJsogKwgnZL0gEb3tPj54azUo6ekNTuRryNcwIQ/bSJo6OhYsniXQg+NVt8O
bBRSW+cL2UKBMTTZveTUYXhgNr1qOlErpsN49Al48vvrPcaBYjovd8T2r0jCvtAFBWBsoN+c+dVk
DgBYt5o5pKHjKRJXkSlGfGoy06tXPs3HjcJz8RC0vr3ZgRFGKTgESbR1bQXLPcYJNDtmrQrmsgJc
ybQIMuY/2TxXb9LMsU9KU5fvDZaxi8QvUOO1E1CgMNdgxuD73ncbnM29gi+q8nYP+66w31z7A7vY
Gqi8p/dAyyn8VtJe4tPYDQjuPE5OO+nPXoIe/FfOz7jPvY8ij3NpIDFp/9HZ2TslLEkiWb+ad2NI
I6Gy8NMf4FvecClFxJGzJejpn9K9tCafidtdKWwWBjffg/XmEr939HibZsF6rcwcGTPuuTIYirV8
OWibicuPfA4rr0yWp/3L58ZLHWR9ZUsW5ciXw3eHyai4HcD1io9VgC9ryvAndddRBBITmJDbWPUg
Hww1KTSULRGk3TLB9gMpOSCFVSVJHAIIsIRJ88MuPoNhCPybqCaxsXVkRE/e2R1L+5xj+fJdtZIG
U0SkBn289hnfjTds4wvE70/QFjlqi7BHMAuidQCUhtKYYV3LYo290hGDUlGFt2zo2MH3rPLlSJji
gGZZOWpPWLfCHLvpPxhNSC71bdICFKEH7aF2SkXzIdjhksjuB6y72zi73j67qQd9hI49Jp3tNJ4Z
npJaolxZym56fKnxmwBDyJD2UKyRW0TyEl1HseRXWcKh9okBm5tHkZ91AJbiVDvkD42H+sUNLjPB
qEJiT4juakw8a36lLnrFTWivx3HfE3ahHMtODR2AEXSoPqcYxy6nf/DRC4LWP4TFLqUOcn586XcX
3+AA+G8kpx4EAMxTlhV1cILbevYb6aq8o+94zrrKtZioiVDpCJqBpPZjKf8M9kGUAg0rf3UtIdbK
N6P3QMsMkICBXPMce8gi9uAebbNgxtj40oqgnPqBwiwHio/T/Si1COB1myEeMoOAeIzuugM51Sd0
Efeil1yoXBHxDgic6hdGn6mOwDcYvtUvk2O/LPO2L4UzTZLgh/Y7i/dsM6PbHF8uYRjPohFMPnUJ
dgkXV3CnNpQL5B7mzN3C0DVa5dcf7T7ELSqLmVwow7stcI3FysczwjhgN84dcT0eoDv4T0OvHOHe
yNvIQqEhanJn/cziBtikcSrDvpC31bj0zG09hDvgGZJUU3BHO8xu8rDE7hRMcU49r0huSdy2ANOv
Lxve3hqV5/GTrurNVfnbWmM2VAU5WpAPWDhzQiOVOoeB5O6UInzdRzzdJRheKcaj0VUG/S89+HvZ
FMs0Ewij6uk3hLeQThI8MLx2ziCF7uXflcn/glm4EtKjmAnJCnoiOmeZdXOjpvOlRSTPf/tIVtpw
Di7iQGxxazplCUMm1VFg/K785yaljvzeVCSSYzrav1FTGM64/Zz6Oa9mh6Tx3L47EfjaB9CdFFDJ
ZGADHb8et8GELw7Imf206eAytUS0AzIwVYhUsj1Z0s04oGYerhUQmpLOs7OFrP5NmcuTuNmD9rQB
0SeHfRh71gwmtr45nKs7BE8Bs2kOa4rHJV4k2WLL+D2UTCYh4ITTLhyEN+S43BF+VM7ib0RSMqQX
/K2OfxxzOei9Uw39XkBEM+42A8uR4ID6sHk04+m3giOwjBzcFz3CDfFp8iSjwNzTXF5GY0q1mQtA
pvew4kaWl5idahVH8vGRhxZj/EfN5bpfK9v6KZmCe4un6fknJV3YkyC/WnLrrYSgzN6BeoydcIlR
eAeu12odNh4pZE0f+C12qqMS8QoCTRmKK9suP9dgECvtLv2nkTWQh0rc7TmeB9t0KJVh9AVsidZ3
zRcive/R2ZDK/6NM5DZqMnAIS4kavUzC+9cHCLENzOFGGbCEWKd9R+uDMPJH0p9+EdhlrjRbzLvh
sinX7+tISyEbwBkC+9M1md4JlZskq8Y7/rFZ0kRl6/+0lyPMZkH9Gcphwk5k+CvIZ5MBDQeCCjHN
B0CPuufkbGnF/5HCJfyp5Y80WK94R4gSznYUMwB/ajHjpDEGyBMIZxHyQJ9VVMly4+mfpSxWgH+Q
gHK4m7ZpPtqXY1yiVHJW4HANv834qekV5QzIjoWtxdwMJhkOgnxaheBoeHUTqOiDIEen9bti4frT
zH80U6rU+60EaPHRAobbrWWMqUkZBC22+lPLydP2cKmAjXYPLlO4zwRoZU54DmQVqX38ou8CY9/q
AuajRdXDabnnjSamN3GYy//w3MjRVO8dnDXDOTE7Z8xR1abnnb5ogx6CjGdKV3aUCA0gnRMIZ+Ls
N/UKN7yJ9Vp142Ofz9U9/2xLlrzfHlOwOq1quNcQhfSE+mVOzYIoFgi3xZ2WQ8DvkqNUR0VmmI//
Y0W9nLJxd89L5luWBHdFLi0G3elxmDCtNDPaOGCKxuiFATGv9b+iwuuyZKuebSuVX0xAR/FUeAyI
uXvAFhxQec+QC2JT6g/FGjMtD+Y08h597px7aqia0f5/gYZQjDFhwI6f1rN38AHSru/b6ll57woS
manKeIYyaN1lpzT/k0qFcjq6zIubT/zB0inBk3S6e3RlllV1yFFrNfv7UeZHEmz11Mau24XbQXXA
/dXebM4rjYQR8zFgAmdQca8T/qgzbDv2i8g3TXtlvf3XicHQA62aJuETKG3kmiXictziNiBnxTN9
/+bRNklIe8DfXWVVEgOOAy9+f8BppVShp67tuJMYyDwMyx3wr7ld/I0slrZ0pLp0fs7wIpKZZRb7
5l8jujqHvOqdzm3atID0Tji2oQApRfc4MVnLl2lnptXV8nqcPilCuQbGeNSteP+dXrqEKg2Qx6sF
CMGHJUzSKXGXIXB6LEJeHRd/wLocl8DcqGVY5CSehJJYvxRm3jIFYXKJ8C03OgrDlRw4t+D4vKmL
ome0QiGg3MNNpzu8Sv63oBRwCmdkUGdTZ6Sy5ZlxpNga1ZP/cQvZ0UyMTcvf8t3fewtaunRV+Ndt
AbDvf+TOh8Od8wRH+zflOBvrs5ERUTrHtbDR5wS8E8skn5n84AaAQpRnZM9nkBn+gCyTiFzxahID
WbSXJq9/Itj/E0reTA9W03GSYiLKVyu8HPPbfZ2fejVQe4Jlazhq4VXRpOjBR5ErCAW+3jWISV1M
OEUSWaG4rhQfXAzqdlltUxjfCpHAChmIUHbNfifgCKq3chZEEoEsMCnsUagic6kC5wa79z6Jpv4X
UajzKYnMdw4pWYIyHnWoZun9qEBDsKqQnhzqXWdywbXD6oW5rUIe/aAYXapPn2PdVEQGDRRwpw0s
NfWj23BsYZAznO6hv6jSizWmnTQ+YJr816kGey+aE19gOrgKTnKnR/Uz3O1KTYp3V5G+FYS0Kqxf
XiUQ2fOtnZhhDV2HdP3YrLSkHU7LqtfsGGXXv6hBhj+D2KuUiBRE5LxksI/ZpkAfajhocLikzMB2
Tv1QeEc+poaPMrvz+9DNUwwYw7w6OX8YlPgwSml/UmtkGhkHsZc8WMZjgEn1CmMVDSv8RDFtWHdg
eM73EscuDs498RXY2WW8v1vBAyGuLNPEWIniDWvUkC3xr8ftTmbP9aXrcam5RwZFc12CaRmGWAwM
OSaguM7TH/DDUG5Pi2K2oN/c/A6Jvz36zzaKEaLHCnR7Wgl1cQHLEE22pzv8WPpZar0DSLbCf9Jw
dj4iQpdQipB9WSqmYmF0d1a/HyhO1+++Q+dH8VosO57hEmtqgYfQMcXesJJoSKmC4GcumUN2jaPl
/liAiuciGHvHm/I7JhzambMu/6DsCjYHE7wqHzzBT4AhR5VUlfuZLiDGgJdEHdm1qQxpdM2l+3td
d0jW5uhGi47lcFJLwdqseKW9t2mO+3kAjZXbPCrhRHQ9qQBPgUUpo0sgihlVPJXds4TZiZOvRRbf
HMVAhTrJslm2NxEOym/qANlzWD6l9oMZbMOkFJ+CYvxCrnSxw15aRddHELuyryRIpxPv1x29SCLt
yU02vcPZ96T38rPMNp/z8CsaPwc1jO1VUWgwzNk6wKEAz3aF5ooR/TJXVXtaRdhLmdruAGU7E5XD
vAzSt3HWNyENaJNbvVOmzjf5fvskBr0T89NxlzKsfEn5+PUqdmUBNVphO0jOUhqVBjo+Rbl2IyIa
KPCxDgeRD439T2TEw2stlT28OG0FxtGc/WAS1IepxyQ3qGE7gE0aqNw5fNH/jshA9dl1bQveLWAX
S+tPHI41jh/b841irc6x6GWYaOzOFdXXgQhES9bjaAC8F/J/kawC9iJPjZ43dG/GYnNhD27YRvqB
ezc2e1TCL1tdAJI1kUkRo4xXlA56XTIseFGwNkwRnh/1BQt2zNP+9QtUGGBAgcwgukkwfVPoPgCg
4o+dlAmtivr27jJc0XP67ydFbXAtQlCUiL5yer3LuOw/MLDAkZ/CVKPeDcNdhkPUT6cxvwDEs0Xr
HNi1ZrUcAnoI1gC6/T2usbKN9WQtZlNGsq9AMHLASLtVyK87e7JoV2zv/wfhWYmI2TGb6GmLtIue
F/0i1Z+b5TREjDHPEtWEuabkSN4wRPQz3ZcHY2ewACrj+DZvAN+grGeY/S5jGzrSgHOZgwAh+Kj+
nERcxW9rqKmUVi3hUzscPoFGHQRhuBxQw7Mfbx+4G1vhZlgjewy3/jCPbz8SZQo5LPhkvMcUzvWA
pQaRY3lM11xnE7gjBxvRK4CPeXKAzdSG4+Cg08CS1/56nUYfMvtWCNmVQR9CZjCjdCIfHh5Nlc0A
d1rrdjdMSft0wjuWarLbLcbVaj0n+rEUnu2HCbIhOOq8FmCCsYKS6MnmwdmxhPchg+9GhBfw9JrI
I47f5Lc+WQucAIjXA4Sk8oVJ2gfsgBI1axmq46tGuGabPbvmXs58tfIjxJq0GSJ2R7roQef8FsNC
Bq7ak4jZh/YbGG9sckUH9LU6X/0XW9kojVUnfEA02mEwgDi94NFtBr6qKJ9LqKTAWZDcMvMzZXl7
LSarT0Wt4mslpeMA3nLHAl8b+fzp6gyW4OgEMlWEu3Rr8sLNEPYmbC137HWa/57Eg/+vtW3oEoeZ
KXeKTEMHhXc/n9g0a8m8dfiA5TN0gpt9CYKMdAsZsJ4MYS88Tna9ZwvDqQ/MDmcWTZZZl/6gdiUz
tcNbQ7+MPJX9Ceej0SO6vp1o/64RWkkVIE6wO0+whS9M9oeJU3DTEx12DrgsZ6ZjAV50z68ggbih
7gD2X2C2bireV5E8yCdC40K1SV/5Go3AHvR/zs9zWuLIe2vapTyk7zwpeI2q4beYmZSeSghLsxe0
Ewk5qyBm7BruA3PyMDoZKvrg343kcgtOILZ5sXQiklKc7+9dy8fnG8xp38mAggsAIwR/bqn0IurL
7fFPJeSpBwlpNlHN+SJw+fN1zz+yBKj1MQzGYdUfh1ss4FS57bUbe8Q7/xdXrPYNecfyLuchEWvO
3baggjgZJ1b4lS3dKBGsV2HHCGVoGkdsKcL8kc4DIEK8lsgejZeLUnkuamMPEZggU+N6LCofc96j
PMj89sFeQw30Wo3eBTY/dpr5NFJ6BLwTSu2Va+7P4qUxzL+4eBAnc6wQEC7Iumi7go+sGptQKDh5
NsHHyEQWGoxjTqWlGKwQnGyTzggB4I/tI793wsdzmpe4g0ahJQ7WlzwDMtsZz18Vz1EP9YYndRT9
1KfV4NLvlqgceNZy2JfKmfZjlth1w5Y58JKrpNqrVMJXY2Elh1gfrWsK5QZPzZ7GStlQA3zcEdyi
o8eXTEtvdwGfJiSt5aNyNli3Sd/3Iso5Er4RNK9xTkcFVqAmhsYlPPSoDZTGjWppwnmF3o7Q0f8U
1A9QnzfzfIxszdU4pbwsqy0+WU45l1wYJoYzSE1U3Rbzc9usMJBrNJjFg8yvbnzbHh5KVe7ZuMyv
25mygSdDati8VABbEH1i2A+kgOp72aVGVPgipNBKkW7aLAemR623XsjJ0sCNv1sItNhpUV9qscJG
1F6+5h7Outdcpccwg4IwyUJLFj9R2bOYYf2JzGQOHJIJYZUcsT9mbhhugcx34TQ4nbPkLkaMSgSk
S9TUvXafqf8OTxiTEUOC0Osh4vpkYoVME521rN9RfGZ0lpC2xfvutQ87WJdd6QAawSmN/V/sehXH
DgS9oanSdJaUlfAbbMOqaPs+pWiDrkhfV6a3Gg9twVw8TCCzIRa8eb1KiSeNgr5HJo9cLbP8brJ2
tv3ZoIOHXdTITMBwgvH2u4W9qSfW9W3uVBVRBOvxcMwYHugIYpHiqzzXMCZlsfghqraLiK/XgP83
IAe3VYY/AvQh2yfxUvslhZV3/jLP7u15UI3hFJXWmhndgM+U90GzPlSvdkqVCJ/+5LAZfXR7+nf4
lGvQGpkN1kLYXoOtxSgPQEC3xFgKA0v7qCp8nvefG2gcsIhCtu91mwmanT5bP5k3+gubczCOZ8VA
tCjh0JTvNBNekXgcjE5anhTEQBagvufzRbw0RWslositOslQhd1PzzFN1dkQ/mC5j0WnDzuSrgbS
dUFLSofPuJOQOIBM5T1l4anSjk0WcSjJKdFkMqx/UuLKL0vOgfEGbb63bz2bnySLMZCDGgyGrRwx
+r0CHMvvfZipmTs6r4KwhGEUJBLDy9HK7yIrLg5SZmGtqS5MHVDQk4Dq8jCOvCMr5WqPp68jUWfb
EwnhNKSh5uyYlpKr0kcffWclzwYImWy7QNRiWcp51DmSR9l+UaQBZNbf5R/D6tqmx8qHcORrIMMZ
XOvbV0kWhXue9dS4kZHcvLBxR8Kz17QmUddVQjy7RCmb5PpZEG9AZ6i3zf97vMIsediPCbZA0Osc
4GYitlTY8JpBCgC5YTQtzVdzHANNk2I0ilW9kz2f6Gtcp3mFqCjNlh2BQqqBw9mDbVRAI9IS6QnA
YRzhYg0i/f4XFsVe93KnWwNaC9c1wTO0IBBb2NOl4hwdmpYMeYJpD9TH/Pj7kPfoU7WyeUQKj+XS
q0jPmv7uNj7s7S56Tm7gocD5Vodn13cqMAdBG2CxYk9PaCYROHx2nq+iVyViU7+mUzu4CgOeazD1
O1Oaa3AXhLKBfUnEO6TzwwnYjOwZayKCSRSEmTEzo7Prjt9N/nSW4EOkEOg2gViuVxyR6Ag5rqpj
UlPWV2545rhdhNNx/ufEMf+7nzW+GKZyenwgSzxZyMHxHFXIYROvDFdAZgb5cdsi2reFptgDXbw/
WqMCuIoBe9+idyBEfArQkfFh0eqwkuvvFiAVJoiGBK8MQxP5ajeiEoEj8ekLOT7pDHkUx1AMBEJh
LIQJLVkx6iPG1QQheNAqmwfBoDEWRqZt2kX7UKlwFhSUoCxu5/TxSv0h7k0dRih8zQixuuPrLiwj
W4ZDAgKl5gS8m7K+uBFNl84w0TI29O7h/2Dm/dmtuOyalU57GRKSfluraittklu48lWxhinCC+Y3
x7igZVmU7JJ+I/eR7C6SFzy7+j04NkYYJ4pT8denoDHbbBifssqfqrWoM9wbTiE/m5ALc22zNd1m
of+JOBUgcbHphwJxEbH3tFjeemunT13PGFkQ3s4HA9v9+OpkvxbC+iyJRdELlWoLhsr6TuyXTON+
Ze9E7Qee1QB5vJPq+U5FJ0bPu4LXIhDaEdWr3j24IGd1FyAZQ9pS7L0yLec3EFuP4G2WAgQ/jifo
T7npq/pwiwaBEDGChJnjRMeDZNBbI6Dpn+W7s60Zbf84IlB+SHV2kRXU42DtYzWoqTRSaT0N7gT4
hB94rQOBWoCeiWxbeWddhVV58ioXK2fchf5X6ygInqznJpmJDYbWHm52GFIdfYtcOGZPqh/iMGoo
BteoLSWxIOXc33wtxOUZcUGmy6TUgZC69PuvFrIbq58xqWjUq1a17W61Aod904dDe1bG1jZyeJcp
VLK/Nh+LJ806ePAVuhGG4q8fyA9qkJnJsfi3YVPSF0GQeRX9WazG2UgOBfu4znXHnEsFwj+TCEAv
5QB87BvRvvZMXLZgxLH2al5gGtSDzWYyopeQzHovp7epJ/Xyr40Rq6XXi3ap+b3RgYcEdtKT1gD2
cVmE3MMqzTYFjULpXIJi/rhEyTCTJIR4JRgWilCP9qYp+bNbvMLClTqXjDRY10yy9VKNYnHyWkx8
v8Fqc/v4ybCtT76eTTkxRv22QgGURP0rjHoeN+qBWZmFNuftdUc50fn6OB4VbDeZ8HADQzjW1eK1
5U1cao109BwJonsTrr9JZvumFB9pp1dvyQJumOqddYYkw3hf18pmfAtuk5DgmiWBrGY1UJXhK4I5
y0vyRXDEgJZe8FDzt77DKaS5KREV1NRXp54EqIC24JnYKbsH82ShC3LHgHwsxmWHKap+g6nxvZGe
ekc7XWjLtyfq1MTZz2qrtj8ryfcVCMtVk2UI9vVxOp3JO+PwXjOKeXkJWsKkVgQeUt07It7awQ5N
8jqvoHKaCsdRD9+O46c99UB12l8yK694JIDiQ9K465bPtlaIslQ8Ny6LVSWIk8ZrpDzvwBv3FhWl
0SON4myL//C7fMGdbxu9eK0lObQ2MmpOQVMYOcoCHrLesEqezijk1zbhZb9jk4SOIXA0gHb2tJdf
MP+eoRuN70yklbdOOeKNmqQk4jqJ0YcAb9llLpcVwc31z3En2/PK/HOdD6h/PpqrF1CBJUEEh+5a
wghYylOII8RVcPshO5EszO2MJNm+44AHWli3HKgwkheihCi/tNCmHOv2OkgiE4z6//CfYrH1HKHL
0Wi+TWT9ketK0OZ/E2J2ftzQzyMnRyIDpJW0tSvtYoSTeQmTloag9/aoAfk1qtg4TjBnzBfKyiit
/itFzUdhRV7Wgnw9xgF8Amw9T3IdJ/0Y2zU4EkBhsYAf1dtCRIdEmthloyRxLZeJGXqALoz8Jlw/
+ADqLTkZ/R59XKPF6Z32XEtsE1/3jRYt6xUSJ0gKPYRmdD+l8rZcyh0QfkrVtGZTJTqDra0m2u1F
n+SnW73Jg7AuGIj5nzLjT1tLyCLCvL/mq0FYYLbe+GJiBqvupmWXlWAWf3TX+IxTPMWqWudp6tET
t1Ny934Uzgmczw3h+aD92tLUCmJSaMfyxaIWXnVEQxIPG3CjgJV92cYJnpeEoKjNjnNnnEZXmVJ+
8fuDkPhsfoXgMnij0tN96nSSu8SaX5aGLsEWyW+pGtbSaZw+x/S+La+LKtFvzhxIhVGptGzzMrWI
jiyQkbo30OLXNabb72vGz88D1Pn1tRY1hraOgPeuw+O1NyAq3GZHFyW6GrUgjvWEQ7+UcqrqXD6i
oCllTkQJnLP6wx46nGiM0pFzwolorWOkTrc8DafYuSKOYX61CySuhhS1pSFnEXH9pgNZWN6VT6IA
HPmaWnLN5DG/27SrtQm/Y+KB2qTpBoYE9D544HKBPxEvnJg7A7daK+6BNRAWBWoGtUT95ppNcbD/
0mg3HsOa7JKrbd/B+JHoBSWU7vsh81uKzeEHysFDkfdG4QwL7v1X1A7zUE+q2lIWH4d7JzYDqO+u
xatkyGYk67c8lcHzTXjlPttuLk5LSFsNBajQf/rC6CEBWYnQv/VRKxPNAarxjz4l2uK1jPx7SHYS
711tvIfYQ9TRCS0+lLlDFHhI2fQ0+pJAtlur7i4WaFbzXUPF2UfW2HIn0LPGLjOB+MvSnoJFnOnE
YhM3j9GL6uXek2ZHij4tWeoeJ0VH+2ngvC1/NaKiBIo+hlPQAOoetK21Y2FZs1bBcMsn0dOwO4QL
z45a9T112HgqyboOm4kDD9OZCmCoy7GagjyIrzGrqaH5a5vOw1nCWh4tP7b+NliMobUi8IIBtr1N
Fu2PBn7+RRU3oedi65O+OYFM8xulNqYojfB7BS9QQwW0z8QLO3qh0yEgz+LElBW+tqQguqt0E7Vt
BrXe4G/YkedLhEgrIes/BGEmcLYx6zcLvorIWVxJ5mcWN3kURTr9BynLKm6bLeyCCuw8x0NFcyAa
5ejVF9rTrBJNGk8X4Bcdg76ic4zQHVUN0919djcisvERgxLCFCnpm2NXLfYLannywwxaX5cM7nRT
sd39Hklqt6DzUAsTQ4wWUSedBWzpdZlhfCFwgrdZxAxo/f57WNYmtE2wum5CStBCQc4W9kN7me/G
cOq0uO/FChvw2RTN/Eji9/byw1dkYklR3jjarzO4zuN5nUJzWVfX3u+SBgMSuZth67/ftjzM0GV7
82JJ2khyY2IrPGMTLZr1nWJBAfJdeOrXwfsKQLSH14pqiA94huB3Te/IUvFysth8atzv7G3sWko2
5mJB9FbeyScP+gzx2IvS6VLAnAzn7yVVTjyM0xUA2ygFUTFgbyy4+NeFRfZj+IdAaUakesnnr7dm
IACfmz27RuY81pBWQungojOeflHQJY/UcObzpgPx9aHIIWvYrVL+XaqK4mnKTxH/JQGBdHtF21cf
HNOQbaeWxAInUm++btwQDzwUGFRL3PnWrCBmfssMy1u1Jc0UthPQENFYpxMS0FkGyGFDai1nxQ7G
aDAaOxJb+nFDfXh4AfWE1MPBYYsT2Ld5lLfC1cOIbwYhWJRsPSYfWgB1gy6OLEbZ1pq3q8qIH+yi
JKCqaMgwyxB7scKrU+RKjoY04WjNjRLFE8OF+T6b3oZCJwsEIUVZioZDcvPp+xC0DXJ3dfuoFBZL
y9rqo5X9QY5f3bgCcHj+H94BB1HM06BdMX1Kzo3Xn/WkAvPiPUouQk0Jt1XqbMBeTpjmknyTa0b8
YpOl/lpypRcr98kAz1Dv1Lpp+JedrM2oI0sFZGHHwdUgtsDC9LoUjfl6ceLmTtAUbIZeDA0BJWs5
I6h+JJAbRO1LmIcVrMHJifcnt/UfZ9hOexCCZ/v425HDCfov0gJ+B123UhjBqQuwyNWoBMG5O8Id
ddJAH5kr3ocXSDkU7x9/dYaCEqvP4UTArEUsLVRUAz/T/q06xVUoelFlIElkmqLneNj7+hdYiskM
RF7+YVkfnbdfMBhOSe505WA6Ia9Brg4iY29pKc6BKaUqJYOnYIGXlQdTqOrt/arZeS1mWLVunWIj
LC2fznlP9FLqvHgfbwb11DIEmOL+OPCplf/PQFZHHXiAa6Qq4+jfQD7YQEqPyeQgRQhRjNRY1YzS
HvphCMjFQz+n2YOIdtkUU1cQjDiFc42c8jqHcxnJ4kAA0M4odqcjtr4c8x+vkytoumW6qluFhuO0
VpgCxxLbVxM7sn3H4Jj+YVG4OwWDT8hA+iNYdyngJbMQojWFlDYeY/TWloRmU5u2DEB7XsbzWHBM
HlgQbuUHGLVPXggu4vAF/N3ixcowa0r1Kb9//V9DlnwZg45AeciGl1Jn/8TCwQRdrjCqpzKwlLoO
LHy3yK/yjYyNfU6zVkyaI1NOtPXGMG9fYzoPaY5qhppHjtgJXiPq+Dmx+z+QszD/ytuFkFqJ6mho
t4OMMfzMqp13yLpVTZF2+uS3Wfn2DUwyCKoTUWD5plSUBEzndg5NFBF5cqdve1df/Oq7NZb7lhzh
AQmMyjvqm9OVqyyapJg3PZ2a+LMtNx+DFUfPkRmLNjLznQ7KAFg5igEtFuQOk/wI1HlolLpAZ4UL
YNVBAVTBI8uQ75F1R08KAonFxQ7LZkwM99bJyZfLfu9oLMHwnQ8w47G0aLMLVW+18r18ZNS3k9EM
sU/WcYs5ZZei87zCipdYWmxnnQyO+Dv/rTbGONHE4WDas+XDDgwE3hyyzfqlkoxzOLkdIiGdHEqx
KDPyV4PJQXAhOEhvvgcn7WqbXeOyCBEo0hVs3AZEayJj+G1MP6M+omvpyEBJPYYDExANu1wxeEzn
JGcOAdAZU9SduODrZ2dyPa/LwAlruquA6yhpb+nUPQP0CZWdKPWjVrRgj7cyc+EdahTs9ZA3dtco
iPXNBmyHou5Qvuk9GjTTxuIifoiHmKXabHBVsllWm5Y8YEmLjFHuwHwpBhnPSgzcjbZ50VfPo4Hl
UlbVCYTi7I//pZxDus4WoSkzDiePXKZMxOl6dclrbmmTe4buUDt86Ady8y4BkGFgSs6l6CKTLzPL
eJbxAYIBDGPXEAUAqe9oVXZFD/KPdCKpY6NHIWulBhtl1/meAJ0e1mljKShtrFgXWVn4R9vY3D0Z
ZHj5phoJZWYFes6Z68J8VsyMWy/w5BXdMTdBe4jax3HKt4nN1Tqz7W1LBqjfigKZ4OaLjGrQf6jG
MFcTJxLLUkYryCwZH6xzMovUDLJCQESTsyRq/ERg0dBwwLv/FJPdb1pGqsUyWjE0c++JERabSqNO
PN3Z4LZjBZiiprTfsHUe+DssAM1ZSIyabKAenTvny1VmgpzhzP3DysDhoBo2cU8kLc+zgCna6zwg
u+iHL/eyrjisrlkz1pIaPMXYP4gEFIqJoAL6hFSck01csKvUMrsvHgHsnY3FZpXn1+TckQV4ltoZ
XHYso/dJPt5m4BJDW0kzPb7XzFeBFJpl3fr3rlPtT/brz0aySOE4HAXVFcsXC4SjkOvn5MaaDGvK
bXaayvASTGcl/JKSik0ASFqxaJqlPrLuJ3ciZsDjNiisDkx/ZzRblvkzf0am/wsl5AaUUi1pX3xM
rwexuSSstrEo3Xz6deBuHadWbmdUj5IuV2AMTXDIvIYgTiHnhPtYtdbTYm4tHmzDM4bn/pJTT5yd
a/dK7SFT6amD/x/kfSW+dhnBFZmc01BadJ4KPi5LV4g9KTiI5VLmj6cBz2QNhJHQqx/aPULjM27B
stmlC66mvw88riP/8dSmdh4uQjOHv3R5nfEPJeSrsseld2IBvvWwkRLV7WMoA3m+phDVqmZojWay
dJ4Un4sKy4R3z2zyaNvAIev3p/xPGwYEtn2yyIqkxjUf2j52+lfVh8j0A/J9tjLFJrK7qvgIuHz2
5WOh/WmEMwcC1OMzSSkbaa8eHoJ0I7z5D6o5L69uOD72az1bPPD1sUzVKuxeZaf9Kfuxn0Tnu4r4
UuRcg6Ip1V+Tlo7W/Aw+0STH68GXheK1/PW9G2sfE0xAInVrW66xrO5lY8pqsPRR3g1JtnK5fdDf
pRWcWTJqbdHVt/61DB0Zm/zQyk8A/u2FzIoavzZ/zP7DG/2GrbbkCWVCaNGe+VIWW9aD+YPbm3K/
BswsnY8yrDnYqlMxtGq4eUcCXQUby3GfmNeawj3TVa/BHiSUJacDggvW7HKEd8wiDqKDm2aTJB/Q
Nm7QLmUtDWWoFmVQiFNHkI+XCkIX6B6oEaPkrcWIQs9UemPngS7dSdoBv2g7WeN4JHl2JaQc0YJo
n1lJVb1c+vPnmJi+VwreRR/yOXPO+/twSp/W0hMMPbI7tMrCZRx1yITVlYDYR8szH+JOg15aQ5OJ
P/HzYdgA0/9evCBaNNXrVXIlSSuWH34BPAJMOzLE+I8z5S+fWnDpShKqXhpxxcOPeW2yYgnis3Sk
t/EB8OaU2yvaLWMIyb0rqKyFr8JhrGImQLEtmdHy3tG0PlmKRW6FwNVBKIzeGtnikPE20Eid1vn7
9itc/vI1o+a4aFJ92T64JdXZE3qO7GO8yRgQ8utBHWvItMxTuMtMdcmfAoGT5wRq44lsyk1zLJpX
fVkBSIH5UjQzKh7h4ffkZlVEb27cgJIO+zu201I6B8bUDAaAakS/Hsc3Q02YPmgOuIvWQHTKqNO+
de062Bw+5KS+0sU/T1nlU4QeNZCRNI61YMzCHn5423R9rI74Y7X5degBch3wQwqTXlyPXWOxB8Vw
MJSAFbBM1HKW2c/N7XBBcnIkHuMD8ry8hIgr15Mzb67kMuyKK9kWGfyDhBEBUsm5CbONmjOW8Hbl
SzSBgt0Iq33Qyp5liAUNoBx5/KZmUVgKli/7cfYupZZ2fiwo6UbW5lSOows1niLfkfALf83hfYlQ
GXgs8UKbQEBTT03+ceKnq3yloA5nIiEpq5oqvKU4Q/nlloq3z5dITSVl41lvTe3ZOX2Eqij/ziEb
rBmCA6WvGLrCZ7ZFHdVU3QgLspZCKuNlg3q7XXnnIf9oCCpa1vk0OJP1Uvy+PlwpJmt0HKn9BnJP
3bE9ipUc2fc2zP8qwjzLdnZ80h1aFJ/CRsyCfqs9okX2Quk+mq9uKMMabS6atN3dLPWDR3kav7qA
Zhf6j41I57yKkij3w+1WicZYGDJgzPlBBWDVodfKwd0nFn8vqTXN0ZpgzAYZFXKuN9GMdc+b1GBN
BQYeBuwPVibk+yDkSX9dUzR8VUb5gmGMx47f1XtUcf+IOpM4TQPE6BV55UY5RagxTuZwqz6ys603
nh9EDw4IGPK8CZPT0p4059Rxj8pLU3QDg7zrbv2xtqbiSiTk4Tf587gjjVcYNAizkvpHHHGePhvJ
e33K/vwNhZszo69IyPzhm6jI5a8tRZ1epgY670WsjzLBf5L0vmJb2u/2d5QmGfTeALMj+Njmv9tF
ptCTPgtKdEFcj61ckTPzwgV013eIlwId0kuZY5pTkYUvnzvDojTdQdZgS38JBpIXrLaNd+UMe3T/
4S5z7Z9VDOJLVpnnKDJuM+MnAfmfD+sTxgNWpnNHbAxJo/FyiGrq4vsF2l8L0h1c98PGlJEOy/CO
ZKgRFnnxr7OI0wGVBf542x7VgmWsMIt0z8b9S/Mkw2ZrylxjqpEGObHgUbQIz5fQHTbKSkoEv2n0
oIOH7yv8jMFwUELqyEF+ehCfvIbdvDd5OLfdWhW14WT0tUS6CHxqerm+AN/2xcz2zaVVE19q7btc
WZZ5/nomt8AbUlotpBHDWftuc1dPVTR6I9yrUMNIPCwI74MHmJLH06n5XOWt8f12KArHKP/ah+pj
izBcBYS3dzx3nyKiTAitizmbbYj6K1KbWNXLNt3u7xWjEaD/yeaDQwB8GCMpcIFLNkCSzViu+ALd
jrkkka3v6oHB7RgYUSdYsmlAmqo/ntooiouhsWlMZUdR8p0fegikONKWyn3nzDRxSp8Xx921ohFr
NiKkhygB4qF7zWAFRTFCgQ3bzbjCePQaqL5PW7xxOl18jaoSSDiZnO308op/hkoiKOtNj2ypugxO
Mq+ZeCEN4hXyQyGqkkfpWkfB2Mv8+M03WiESpyDL4ELrTicQQogOfZC31BBx0rS6oyOlQdllOsaA
TlzPLByRKwZp0ihxXmx2Z66d/VeXIlH4iV1GndRSgQQhZIeVaJcEjnIuWTprPndOMJ9ZizCnXSMi
F4tyj/NA/cYKps7oMLQvGnYGe60dBs3FYtMmJw5qJxFEPD9eY+enfsCOrbVoBD5sZOp4bEe2j3mS
/SfAqpetnlZrVu+B4KIz2owjB+AKlb5T4xpgn8Ke6DascYfvVBcpmGbxH98U22uLcQcVZA5d5OAz
p+WZaL1edTOd+7tM4hTgzCmK1XxuAnyMH1sYUY+0eg4A6ezBPmtJdyHDO3hMvRwqfVlKzhDHw+ar
PTQDAt0ZDtYStxXoXTcECrpABu9mdohSFyQgNYG9IpoSHpKF6jXGCim3GO00mVBCThskEO31GWkw
hl+OwHaC3Mvs1AL5kpjJZCZGCMV7VohwP8xwtnZu9T4z3B81auVy7UeJM6hZ+IB6K4KICckv10SF
grRoQ3W2S4N2Q6gIFAjZ9FNvostyOoCAUdD8OsObvN3kXGgmo+VIMe4LLYeSEiMNiAj+rZAcW1W3
aMJTFnkVsMqYh/NwvKdDi7/Is+d03v7szcqzRtLRN4Be2rxRE8z/qX8taDkpgPKULIJK4YuV+F2X
5uIRBUGueyTmjhhFUi9sf1+gTEGaZpZ04Eq4AvC7EL+mo10WKF4yb8WE2gCdzytHZPXBangYPPtY
tnxFPUdMSnZh/dq2VJID0Gwr7E75fcam1tcIiECrD9vRT7/sCxOtPXbiwWNg9ktiS3qLqC5LcHwb
8J7Kjb7iyit+ZsZ0JmjRGwDMfW0z+PyPrZ7tF/PRpQ3r7sCCuk7uMktoLE0qsZJuVuGAgDMTTGA0
lFfuIrDTrPMRxtvTgFscXyHLovBssPqMizVlRzMDTjaBAl79zLKj7d1TNdjpOnRxzjPS2P2/hi38
XFZj2bfO5UBkVRK1b9wPciilQVisOTPf2ldz3Jl3sUXQuywjbCww1LLDHXJoFpDdcwJFLwL62tTD
/1RRhkNcpKlkUKm1n2LKbuTnzvaZ9yz281cqpqUxOunY+VAWIk3vEPjlPkWIxSBO7R97o7Fqkn8g
1SmQ6nGALEgzeaIyVBqxhhDP8yZps+Jhy2r1p/xV8HsF9np+b1WfZjWh/QLSCGXPOTUKTgFR7LgZ
Jc+GnMThl3brgJ2fQoLHjGAlUonnCUhkDpVsYMwHv+D5qgoE26gWvYbJvuzyRdhZdvRgON0Op+TG
5DAkOeqeeLXMMv2k1HuluHE7dUue4HQvfE+024zRB9FNqdIdd0KN2ZnTOXl3GLdR3LlhNVsg76EZ
XvCrK2ULxoUWFvERn/mg2bRWkw2MxrDy26MlTov0G5IweQ7jr+bwhRP/DI2iJkUbH/8kMfaB0GKF
VEdZ5RsRg9UW91uik/9klEW6L0qWZ/+4WqmaYKooSJzKFtjyu0Yu1e7MbzOz6VyNggVWkocP4zsy
nf58rCiTjgiSTAMrtLF1Npt3c5rUTVeff996B+hyygPeq4828vTa1shQ/KHeFcmM92yFrUexW0ai
ikli5+4Y77yhKVkmILg+PySx0XG8HMq8G/SCES7sXXjw7WWxq1nuzbKYwacKJeLF3Eq2kNGDE0lI
gP1Ovp49E5L3vPC8F7OWpTlN7qUjelvLIcdZLcuHEOQodkqnhBl1bH+fP8kiZDbrMniJQflWJIpC
pm8u8qgS2rvMLaX1yJvlm8guus5lg/FY7WKq6fh6MKbq5mlkErmE4he/8B+/Adq3s5cAjHL5jOnv
RZdLPmP/oYCDb7ZGZOdoIhQGB59Y8eIw55EzwVLjqkSossL5tlLjXea+aa124tDJsoyexRwik+4M
nx4J/Eu0oZamm8JSfD+IuMy5ZNQT3osVjnWhbAraWJMCu5GsRQdoUm1f6rc4lV2Ms7e7UqalnjRZ
lUOcPsgjyRvirj7SzHdF2pjYnvEyBaRXzvKH0zR/6H5mDGEkQYdko0aNDFAvwE88mOh2lJ5MG7FC
H5sRp7fdFVng6QrX8MM0oQekivI+ZlrGVsQZn7s8PCQSGzFIXSs+vtEVPz5SBPhjAojXNnbCJf0N
+OoI0hfihULy6ZLnEjrD4Jz3X0RLsmTqtmkG5X8ec0Ulzuw8MlHumGH05b0EDJPOHOPeAx9W+kug
voLVLZCgrdo0iTlybcll31GsuEwwA+tF89fdOxDm/TfFH6QHs8eNmhR3s0bGZWpcKe/15k0F/Vpg
r5fc2PUgMjjCIEQZs11uNDKiYiiKEGcwAvV9Ty11SSz0utrwZOnlNzSy1QfTN6Nlfy9dSfmkdDCP
MFA97Azq+jL0PhCXI4v1zh2o+onSik0qKTQ3/hZH+z3wU7+4gP2y3qNrBcr+4CU1OugsKmGsq9WM
pDl/lcT0nlEHt4KMFvcgBRfZvz+on7sraSUj/XVyH2bdzgkLG0L6blq0XYTzFTgffcPw7kNlJRNC
U5M4FQi6nWLSZyVp7ioR/3FMLjp9myawuvuAYom/hO6AdzjDaxobypI2qj0X/2yu06DMJDWT2WrB
gBKPcqAV+LpeRo7veGITwIkppBisp0mp7KAgTb1ZsLYAESvL1hFF0ydZqQuYrRtoywSObsLExyJI
QaQaTJq94eiql8b5VoEX+61gtWa6OSuK6HRCxtz36jkCuKNf4aeMl/Q+pphz5ZNhqcK5WpBGDe+q
RgpBGFpk15SPtdBDoaRiY5Y7Pewpr+JDhzMlehqsUHR6oKf68Ja+MkxUVxBtSzgohrW+NzB+8lxx
tUmzg2bR3YAnMNf7vmZuvpwcy1Vq76v6qecUoRlHopCKkig8HiV8i3lDrizx1wI5yKtM8SU3GSq/
7E+PU5VIk3BeCbnge+WfDH+6L2ikSFiGzQhGzenGN4Ahr64CbfJo1KBuJRsPJOGYLPdrXx0Grp1l
I4OIaLALa80Vp4qN42JestCVaUcLnHsDwUL3spNHtG3BLRXbpfyjshQ2dvaKcQePt81X/0sT313n
ouKuCOjGFM5b9dTcgSYUr7XAr6NKTfejRgrbs3DmNLf/8c7KM710jilUz5MDvF5/hrPQGZQ6KsVy
UmQ70qyp6Hc4JStJuiyujunO9bv8gJ32yaNO+T955X9sGZZrS5n6h+hMPJ9gAfuvnjHgZM8Eaqud
gQjNWxaaM95IhlpEOorhuxTuBexdDo2KQE690AKd6RwVlx477CYsoAY0dFvAKtFI0OnDweZhwGx8
kSlmBrDe7yn5YjQ0c2/1gdi/wVcOf5eu+A2YfR9LjLAISQhpXFsUfav/s0I0oOU6zCpic7gGuAIe
Ty82YwWi2zJswW+3LWczfrY+S4w9WTqckY6xx3nsruJ+l5uRkpJzdSx1UtdpIa2i0eL5/8E/eChi
Pbi6qTrjKyZ+jOTZew1A86lwS9xD6tINne7cPjUp5YvOru37LKNdeG8IZYKwbEOjekb3abF8iD4W
8baFWwnP/NIoYWUocJV1BGXHrcQuwH1BcoAhGoNz6ww8dm0QpjrGU3GB52blL5MIqyS/wzre3FHn
4rjynZskUmID7WQFrDbob3F2Ej7x3dHEBq8nSA8XXrmX9/wcwD1NV6qyKVTJvLVgC47pP1kFQe99
qrnXVk2pLjdHlrGaYi3S7q6WhTBNrWLfhvINZXcCqbYNOjGONht/m9wuHahWq3E0zFyJmNMQ2ODu
WXa/WYrpCQDnK8ox40ahNJGOox0e0zNrldkuEC5VVCNd8F+R9LRH+lFadIbGQTGfAaAKv9Pnlwdv
lbNzJuPJtHzEuaozd2DR7zynYZj7sHXCGZQj3xPzdIzxnllfy5EkmAiUm+rvvvdavLuUDlbIGXR+
ylnWPidfAhX6lS++nmqKkVgkoPL7iGDFM4ale2WRjo6noSspz3H7ZKHEBPxc0At0akFlD7ZoAYM4
NXDS7TziKzA21ZEhFsSPGk8ioeW2nQxCvX4CkUxf6hZFa6+RVhPwO1mKNFvdex6rGLIapeq33IAx
xXzYDPS9oJhf2gUY/xIc/yogiDnra7pzKmfEnDJh8xmwtFfg9mBYasU9uRfAvpx48QnfKcng3KLv
SLtztuX6429UezRyTx9JtntLNJFeuDsFbcC7BYIAR+63IE4gFf8myHOKyhhIPjAYCCuFg/8symId
DseoLbnKQP8opvV9rE7jty3l4dWjboIbIjyYL0V8Ubdx8USMCEUEhjIbvjMkd5Vqpbjeysn6cnuq
KOjD5C0UVPsYEMBRP9K3Qrfr9gvcNYPAG91h0suJUmQY1ij4E1SYTJ1N2bpV4FW9kpgBGyi7pXwk
zP33zG/QP57yFVFgIiewkpRYgjg9A9aZt6aDpG2Vky1/Vj5hmRZfe9cR4OEM57zufXWnAg1acefE
JTsxQDVWRdyEfBh6Az+YAkO+oAPFQKWSNwQrUGFguQoX1EkGuvixQHGjO65zZhb19Jimoald+0jv
Eu8gkE4Itispk9Z5eYGU4Mpbo3SbHFR8gL/QnPQpPjLeahulCXFuKIXZsI8o5uWvVNLJmTIFUkYn
38y369iIeHQAxczx5CYLLwf5BTnihNcbXGmIyWwEUORYzzMkGaNmpoq1aRGarHj/eb7JEJ4FL37U
wuZjG3I1jwwnkpVVlRsjciooN9EhaZCg1xQS7k5mjZ2aHVUnECBRB9uutXk8ve3xhQfgZgxqRF9+
mp3zjgVB5cMgn6Q6IXt96ufE4LvbUpdQCVOyzPK+7MveJZge4PrCozKatxwNzVx2bMPtgRqa/411
KY2E8VMAHgrgchzqo1fQttVAD+4TVIwU8m1c51ZJ1CB/RwC6ELKNujInP5J5CIhq17TIb6ndyvq/
N6uxgxV+dJW+YX2MjZmiW0SDtzF1L7z97DYkJk+t8y7+xF7W5sIvBzkSaldIk28TtIZ/OtfKCKf3
J2LUh4PCPDjDySGTSFGYqXyQsaU6j+xFU0XqYc8nKwpHYXSTuE+Vwnj0w9n4i0SGjm0wA1DhtEB2
nDyygR8qHkR+cMLoZD2fu8jxA2HA9dsiUxB9lCfae2SA66rsboV7nkx179z0o471oqufMFtv3VtU
GvS7iF9mKQialUBgG/CK4Cl1O9L6ftNAe9ZhQYH4Q8jPjzNY3BS9R1u9MVEV1pGlidjRPH4lMr78
6RXhfAkxoZgbc7A00fKFfBJGCM+zbHqMrQJSZ4JGMIe0yk+XQ/NXxXBFvb+T0T5VrxVPDmRXLqFo
63nitIuVY5TSlEuVaJjHl4hIr4zz+rFDmlsqpKHndO99JggAX8QP6PXEqw3qKAN293lW1jpWGrV/
qlMjLRS58vaOhZbwBrkkeJOEauW6lAihztsn2sWR5bpiYzkfUMMMWESKTGBsAjdas4VcpaSw83L0
iIVKJSKBYgv+PBZC3gcjFnZ9ReWCEt9OaSe3riP3lklOt9psfWvnl9X72h+8DGPTExxnOQKUwfrC
ZaLBNTngFym8iWMxDkI9s1fQ3iDJqq1zbQEyn+MRuHxA/Vm9/gY+FEkfComl1sr8vkQrBepMwKQb
o+9sZ93FuBgZEAjJeDalJrcT8aI1BsLDsar9PKp8pIL8qWl9U4S70Ka8zcfEx99vUhaHCIAmQnnb
Kg/0hsIl8NOKBLKLHK+sUNgLCECcrAz9spM7hB5qU3FwvdZelSWNmAKZ4DkbcQy5c+Mx5lkEzpVO
X4ccW0WR0H+Ejg4yqQkVqKVY0l0wMpskw600qFaWCdsEbaFBM/p8GN2NuJCiLc8oU9jq/jrkQa3A
grqhohUebJvBoIpvzOzyEQCm6n12gn8b/WZDEixculI1zhITfNvX2ovZrcPRQxG3fpFKqm4BRHzc
buDqghSX4tZVFN9iDHyCcuiAatafdf4LNI4yiLl34Xatk3MA8spXBdHaOHWYZXwtCWX3piYJgPxj
ZjguI3sTP1YZ6vtl7w2Lm7gAoGxGIjS7/0hbNL5FC09lrubH5nhzFh8ntqAIJY4/lZnEu6qoicvn
lsmgEXMgM4cfqJJ3oMKh98PqvZDCwKBUQAccpz1+1VON8v04n8bZcaB9OuvkmvfNOJ2qXuMgZPTg
t+r20ZvgQ4TmRYGELvS5MtqRzmzQFd17/ddqkHtafBQ1EDDIoUgcGx3/DR11rbe4ioF83Pztwqhz
pF/3/NmZubP/4L3mYujvgqJ6B7dQN2bN2KQjPO1H+S6aTAxOb3vsZOoDeyiA1Pc4BTJQvnlRAp70
Jh1723SH4qSGsB95QF4EmFcL4BbHlqtO1WYVipEuqIIemomDKTiLEnGIeH0znx5QquJeLu3O/cTv
z6EfpVUolJkuTqxIgDDDdEtTzLClh3aIAJ1hQXUOJ8prcciA9dy6VEx2uxgtpUfBelQ4WUGiQXX/
xRgImsl1e1SYAomyVX1FP3IhwULAyJB1JD+GO/vWKFu603R8EI/MVzCRKV+CwhCRpkV1BOUCN5Ax
s4RYH8GFhwal97SqVuVy+T0ypeEnntVrLzN0sjB8f3SMbl6ZqnQPHnqdvTN9jT/JzPJk0GIZuE/w
2TL1NcPFdHi3pQLBQ7sMpRrEaJaa/8EcKY35q5ZSi0lA8yN6BOm8vzeojYxa+xAMX0gm71pjOOg8
0m1H3Bm1bhTfh/Ux5z9+98AYzLYaNYZHgP2wUDGXHmKvIFGn+XKQkGmTd6+V3bwAheCCuvNjNqqw
+SfRZkQy3eT6Z7RA5NGaeauHCghM5yFQAxqipN1WsO3ISnmF4En6oDjPncMpZzZILn2x6bTPLAN4
30DGYBWagZpD/kvt+WsFcbGf8c07/b6IUA2FDfxAhxaSOoWY8q8V0RZ1oUzWIj45eDah/EQBWyI3
9ja+TQHE/umcxWGYpLQN9vl6muHCpT4a0wQmBo48PiK1kJueTuztJq697mZRjWxc+HNYgR4T41RM
LHwNs2djtyMcuemucrD+Tg0/mOXuffeBGjTjC87q1zpxa2l+hPmTj8B5cm7L652JgDOr8yRHKATb
gcUie7tPV87Flpq+9LYLZ0DgsOdkESOPzQSjuXHJkdkVcQfdcSFZArmXqZmsLQFqlvQFC880HYjf
hu0l1k1Kkhl78yN/HuEz+jtsLN1+1ToM7/nmiKPZtk4uS40NVuQE47xbz3PrdwOegFoPm82QsMoo
uPG3fryyLaqFsaJTVrMTpwQVVJCgbDGXXhWx26Lm7o6r5t4Wd4fHpj/bbgBOxlqxngPtEzOWRcZR
FpGqodPl0jjkdbzFuZWhtfw471SC+YNDVyhz0T2fAOOCsch+wG1kA5QGll0rBZ+ut/DOmxyujSr/
tKVVhSQhyVbEOg+z0XOEMDB13UlxLNVNMgh2b80P/l26B5HnNYINZrx4HrYXa/TxL5NueAvTPcHN
jsy95wvDngLOeZgEDULAmzJnRDukid4rCKAyLTh9uTe11yBhEVeQ/z+DsxlzAcHyP0y6K0HuqWlp
lALZD1hIUp72mlA+dqaL8NKnsbL3ms2/SVMoZOdjyC3axA4soh590XRGZXGj/djZCuucC5HFulI9
pDoW3QDYvVqw7L2KjzyeL+PFX/7RuUZAm0RK7ttmRBv9VKveguUHAVWrzOhL/Y9D/b0aTv4XgI48
E4VTyFBXCGjQSk4Q3g5eC00fX7es9l9gk57sdC1kaGmgaRAi19+a2Oz8eafI8cc3DFtvBDt0O51w
jmRxYvohes8aLT5hzwG95Nj0nRpy8VoS7Bv2ld0KDEnRV8T5lhqRx1dDAg5daFhanc6vqWWmCYdv
o26XPU7yxBGxNA2iopyU1HRn1W1CRUQgGBoB0lqc68faEOsCVGkjwT0pN/spjRAZOACcFBluWHM5
KB40PUallxNAO+tIOpUafdz95O+nsfG0kCEhmMFlg6KjHC3izq6WChjOa8o1ifaYaYEQlaOJK/4w
PvHfLsbActPmbd14iSHHgLQFK8271Bg50rM0/Y3YPe1sE/jKO7EQgl0sWpaECC93pK3BLSsIGhOF
bckPuPx8S8x+r9V591F7FWjQnzx3Ej4K5m9ILG4vnZC0BcW+iV+4cb66UQPm+ysqiAHQ6YVoRPph
xn/IneQQQFS0XEvoYn5FPPkixm5eILMi2TmpSrBgDdVs09XFxSVMXzC5U8pwY1jY8shCyE5OHcTR
RclSIsU2dmouv6UrI7crQmPHz+ffuhfB2Po/y1x5/xcVxn86Zyh5lNd5yD74tX2RBipF3iSCgpCF
odr8HlUmRcHW286EmQ6szp+K5hfv266DHsSbeMUq/NOLIMsCZDXuxU7XTBNVE9dNBGQNGTF5dRcN
V0gWuaPFxcsZ5hRyGsNU3Mlhd7hLt/330/JonwXwG5AowS4Wu3kO4cZ7R1MbxsuSeEhzgl5jIeJl
sbeSS1FkmlP48iUtGyNiav6LpJZk721BEkOn8y7JYbQ8KiVvjq2jj/Vkdbcubq8CSl5KD2wlATn/
Tlv7egqAnPdMoTSbJJ0PBV7ImMsVvXieThiN7XfkYUfB5U+sLSoEJDJLMCU9HPP/uS9dxa2+s7WL
0GZs04Hvfg8RP/33Khwt8ZlO1Bt7bVO8D+yYDqUIlQqQJeP74S9fJTkIOMwpqT84/aDKnyBKBOQG
WeuF9hxT1jEqVWVmG722nVcv6vOIW2eJpiBt0zgZjN/5oke3+B2MwRWN40TbHx6DOM1CrT1pUpY8
dX26J41MdX9F56oVT2oX1k4AgGHX4/3x56oYV8Mc5qkYP4YrRO+K5BgWhggHm7ibLcaCbCbF4C7G
Ay8W1VIto210t63IaAlDAdsV6wGoArhuPnjGE1wfrhc8EkneXLmjUaMZcvZfUtIblboiGcti0jMj
+M/6gzyyPjPAvKz0aqIwP8HGkfpFEd3gCbduP6I1/0H4myCLWj3OgomDjW4Ze4H36FZ8lpKkqzwO
26zHP2LaPIBWq9y4B6VUma/6bPqloE1B2sBPD679WqxRBKfCiVQkF6WnxnQrfWOgLPhTvDjPfpyM
cC+bp1UXzZ3m/uWsX+OG7kvSPEBtTR/XyfdcWROMsn5L50c6Bl6JC4x9EKjXz3JOHVt1ai1EcS9g
o77ohjQsNTZsmk4sJvNzjlrY7rkUHxGhJOeCnb6nW+HgRkwbzreaxhI98QufqCJu7nfyEmNd35RW
cftWduvX3HcFJAO9GxGK3vXjnxN57Tft41qbplwbw78/RtHBfUIroONEWEXAaorFuewpbBUg9xHQ
IneyHmhcdHlGOcD/9iZulVBY1dTGZTJ73gifdHko4ip4P9FwektT2Pavu8AVxh+jJ4S2rNX5g93a
5XmCSDVvu4q/NccDbB7a0Px4OTzpDpp4kIYpzytyQfVOuwr3WXq4qQ6cv68AcI15/Wynk09TsxCi
OKtbvsMwHO0KGZJ+qdQjlxJ/zVarhDcddWhRH/gKbC3MonfC4acdaK1JA7zeiRm5zgQVSJ5WC/u/
+adpOCuT6W17sJ6flyms4PXRAhsx4hd5ZQT1XNkSyKCxX/syWtCnrlsY26hZkXknGogbPfdISIM5
jDtwwrn/zvNMfc/FhbnEnAghRDNeLCe6UJkSOh9+DSRFIMC8izExmlEYs8EEtMyZME7HkWNR86uL
G3JgJLZtucdBny1wxSifC/tThkeOlnC+snzTwQxDhHFXhwazlXpOryKrGVyyEQvoUn0iogmfX6rL
ymHpiu/FPpPbd/BBqrtubIdmQehJv7uGi4D4Q5ObSes5E3i6YY2dR2Gt/E8Ghfq2FxaFOT0umGi9
B3bjjo56081Qs+q9wz8gRfYui84KbrIa2cbODS9b43ts4YZhcgrxKvGcfcsBUbkt9JPa/1jn8bJT
m8kph3L71oMVpBhoibs3Fc9jXV4QSWb5ooIAfiIMYh1FRDKAExuXN6A7erW00HkjFpZIPB06ERYv
x6uC87bn5WuIhgnJWmTIaBDvuRc+pMaa7gwERiKoszqNWPjZLxZGVNFKL5ceWn9REt7Q8+pCeCeW
3trasxjFOmcIFWnBUgQEATtjvIej1v0Nex0xsnBk0I/jxlHzFp2GVqti3WPuLNQLXvqXfMNpTnRz
VYp8WP1v0amD8M2hliSuUNUy29+E7s+45dP7HCL5pxcIOfcAbQGrz2JI5i2ziAIC+1v5EOAROLwu
XzNcqmwIH3392j/q8yST90PSAJfoTzUgkML9y7YnCJBgCHGJMfEoOTVJhhDS4QR3ex9oOTuRps5w
vfJt0haxFVakTgMzK0YNkqAvC7QyS3LKss13LvJcOxRPmNVPo6ecCMhogqIiyjloCoHhKS34/11w
XUIcyXPjX0/jdbc0u1HQVERXkei/Ib5GDaVrmmEpxhP2NRpqU4YbUHaqUa5GLH3K9RzNHaObFu/7
19dRXT9wN/jiWCXShKclbmqZld18puF5j7FIUyzPJboCcY9HvS94GAkJojfGPF3KwH0bZ1Ikje0r
1BIqRG5LTEI9MxkqCkrtTikI67cI9kEGco5EIoklgc7q5qkUU9LpeJdM3XHdWSmxWBYXPRfC4Ake
GRuecpbVpQUVqscXNT3+bpLIBEGr5hHxqfk7q7Jz+f7AIALaGqdfUiFmbE0QcZ8sCxrD/zDXHNAX
MWB5pALJ2cqayyMGHdiwhVdZ/XYLm9qW+rA2xQA05ZBb2TQIaZDD5Fhu/LtARmWivZsWP+ODB0BD
6F4jQYMKZqSjf1qHQxMgdw1NmUg5mI+DqNiIgQfQNXPbHBCvI+8JYLZMGg/VzJzmihxapiRCPkrV
zMbWjWbaJs5UkNTjDXmHZP8PediXJa9GUyK2fQG/D6vP2fUXbYMXDvvJ/wtcpnNDmp5lEPohAI1g
IrF0K7Z4UQvbOTMvNugmfaWQz5seBO26Vg1bZHZybx8Pcwc+93qz7PzeWJB6ZVK8hXIIVtpMn6G0
B2zQSPtlm9GBulnyRQ8oM6AgmZgydRHd5PCm8/FJ/YDIm/942Jh/sMEMR80+mi7tvB6DkEQfD+/r
E5ANSDrRRd+o9sOAkWjTvuT1ZSldagSBQZ3au5o9PheCpsXAxo1UYrLTUh7EWPbIC32pYEApwmn+
MZvpOGHmJroVxOO5ufOE4zVXjURjPdBkf7kyDhv1NGm8UatSz99cE7QvB3+Q2NPLnRIIgKaUD1BG
A0b6kx0M5EOVgSRfU4ai8TehkOlitqQbottbMK4A+kr5+z+Mw+8oB+Dtb2ewnFVr3IRCueFzAnGq
d/0tqTYRvk2KddlAsiAL4v7WcChswxH5lQPobCi/ajb03n15qe2sUoOq14rBIGTrgaEStf4a7o44
myg0D+yVNl+isuFYIr4B9ooKqkLohR9q8oWDYwv/Xb757rc7h1MnOSJAcbX/FfPvWFMFYTGiT2Pa
Ye1x0hF3QC+wcoGVWzyOBMrudzNFg25Hu9B/8wRrFeeI0EYY3Hg8otLkZPNWuxurhgVeBqWI9oUq
LFu9n+aUuh5iYkQFiS6aBhxK7duGsrDgqW4NpOXlHdSb7Z8TjfbVEPd6DcMq0trzxnt6qaXhHze4
tmTPvRvzU/a8qerbY0/hLbCE4iN/Fp3lmG2FssHoQoYkO4FIierNXlgAdIbaFR85OiXuzmdpfRWG
80hMh/5QsXDIVAmtbdYfTSdImjnByWXJ4yYjA04SR2pFnCuUk7ciCDt/SsCW2Q1TubCgBP8gi0Aa
98V8dAJ3AUH06BqKaLyOVuGWpRklDUawA7snvwPi3d1kXZ/vHbHdU6pEhc8x1BetUpBOt0HY+xKa
VvS4VK4DewKenXdLLchvLJMBE4y1SDW70nKKVUXMsdoDURVv3wb1GMrFIj0neTUeKG2hTxpGopVy
Spf9+yltgd4zAkNeQGkJOYVsu+OjR4oYjEWEky8J+4p8KU5vka8R2N2u404jTRy9fm1lyKsPD3KE
ckWHkeHSnSWAOp08YzenTlUZooNQHqBmjYgnVHB8fXhbgs83Zw1voagYVRj2Km4SvlO29oGnJ/UH
IAv3Oa0j0VBFUpRmXhoW8fk3RYuLXPAxEVq5tGWLZVPdDkaC95cxLUZ+jIigk847QRH5Fcip8B24
JMJK7zx0QqSCl6DG2qDza2RBsumBrM12T6vznvOXHERC7FxdsRl2HEMZ78icLWXmHBO6nKbWMI0y
xse3Ch6VglqzRoYb/0r2DnSz7On2q5+3ba+cm382HyAVhmLaK7VMu41hNKQ3ZSplcWkaa1w10OFF
PBpzmiI8b7MSSSa01zhmq+/QvZU5Y0Q/VhTdTyhAUnP1nXhZKrs44DDihRwzDxWuEXV+knSMY+C+
QyqBXmPoNCHp+kDBt1lU6YH0RF9CE8VdJnrquHxQB2880XdGZqho0FHh2fLeJ/OS/l4cuRIh4281
M2KZk31PBS21CyI5tv9lOkIKFzklLqfYZhQRDkMrvGUxHXjjRevFy5DV5qkSV0vyUCK35lK8hVsk
zsXgW3CuyK9SKhu+iQ8dmKqvlOS6PoPqml6XhQ69ROg6QfDyW6F9QlSD1Wv/JvCn0/hevP+20Lcb
+mrpouReMum8cFjiLGaphnylp94rsfyYde/fAozxcSrQFaFZO460AUHeUI0ClLW1Wv3fuAC4fMMb
fe2JwC95VTlPUOeNI7qpmHoZkZ/B72FTnDNDUDZcrMtTdb27TRPnPrA+D/O6TCWgsf41ttG14mA6
hbruCWBUx4r2OOeI1pAAGs5InNe2Nw6kG7t/JsziePfdlj5ONsWci+EyoIGrvKLbuO4JBjbqVyuU
CdADPGnlhhqR0s/B2cIHoENYozppHjKykf/pzLfnJe6H86DJSohgdgkTapdmWmp1RM8NHK6JZnJ0
bO+VWMN4M0imSlhb4kpAGSgU7LfWZTtfsDsQZ9sMJSNgenf+qtcRomacogLZ3yzQwdxhPCUVG37X
ufZMVN2TEZY9+DBZIKRzdklzN5tItdnHdl25wv4JsuJ0I/jci+9XL5E735iE0yPgpwxytmKLqp95
1zK625PvfS6SWMvetV2bkpZ0hA2Jx/AXFWElz98KQKdKSUbBx7pW9wpCkI5+Gt2Tq765kqIL5zau
HimuQPBeSAHEe0ezPER/2CKoa+E63VKXqMw8Bz2u+EFLZYGSnbJYo+PmAyionjYVJj8VjHPHQvKb
XZqnh4df5NFKrt3rSF64Snfk2jj+o9aSgb9w5tpoVpmbuOb6KI390Pf07OxTMwVs1COeVHumJ3v4
Rh8NHzbqEP5ZRzk5tFpHFPWbiG9UNXxXvOiA+VR2iT6ZQgwITimdN1lKG7+OuNEZButJUMQDHoqY
gVaGZ5aROKWo70RdU9igGquuQKHO9rCSKOsyjZf01vTM+9eUxkOiVoRQkChyLzYACfXeC/cPjcTR
cyZwY1f1sAYOY32QiibutcURvlOYBmqHcqa5RYJzKntQjJMiQGeN2ivWjYoG1RCp5RrQqc9VCr8x
XSl6tf9pm1Kw44jg2tLf6TRdkVK6n65EpOt+YZwu4/r+OpOpadMUZUBWZSJeiywH9XUK+fLjgODn
daV+/ItANKt+t78faDvQSIBvqLxZ9RV7Y6HoUuGAzkygXINA2I2rtPeIWBwItq6sOo+DIAqU491P
wLltD/IhEV74wR4COCwJ7zbmUgJXnVdefdPNVrZyzu9teRbplRbw8mgZq+M1spxahJTcFrB/Qnbn
rHZHSvzPMbJ2d/cRGnycDtngIBEQ1mfJlhVnte18TvPXyNf1THtv7ze9j99MPwYd8gM3003jf9Fs
QAvOOPtDJi4/xDWtGlAqtDptovplymu+3NGdScuZoNIT7en3Ijp3noxyKoxMrE0ZF+CDVO/mscGS
FtVZeQxoLZJfw+Ey70Y5A484B1oTCemlP86ZrkUJ4QtUsihb91Wlpm/O7uQm/YSOnjADnKBSL/qz
DupPJmbU5Gx2jN5tnY42LBX0uDxrcn2Iaz4gfIYMLOLotB4rarh0EsiYEy+YLNWMGY6b71+WQQCX
550/KbqXvoIMWjWncsnog+1UEmLhsWv40GP9530AWuhE/NIuge0r4/1d8R3DWmwgd/JOpei8j6Ov
6elx+ZAlWeQOFGo1SWtwke0D/FsH6e//o3KwpA4O9G8rAuanUmzN1nnYQjGAST/3mAy3ggSvzubJ
VVFt0s/pJ/Xk6P+6Icz+7eR4Xw9ZLE6PyO6e/AW8g2nWa0YY1xgRnrrIajOU6P/NEyQ3YFegZZWy
0g0tVNyfkbPaM2SMwZixmB/1R6KWuYYKARVKJjhsLgbNhiM8+1hm6ZtdY/yExWux+/el5OPQssz8
3rLGOiOh4hD0ZGG5YsuF8/5FOePLgFD2TXAWcqvEOsZiCCLWhSUu3wyWfeocTSw/K7gfCByevez0
6NUDJocw9Z79LkgEWuf+D00zWazDHTMDhaIvn2ksAe09ukWcLMfpCNC4ajdjAm8Q1lXSL+4c68fb
o+K1kQDhkHHOycQGZoO/OUPdIgmnqA02X4AHsBFusm0i8bAxLVeukheikXQ38BpFfAEjhXb7JedQ
qNgAANbI27WElQ3LgeUmw3DIlvyQRh1cvUgpOLP9KB9e/bugm9uJbzmRyEp9CLQhOnroUGwEknWi
3RlGp8CBYoSZ/DC3qMjx8oU9BuK5/7//m4sHDxQPZImzposW0MnJeLaMv7jLKBnIFb8R11kBXRoR
6PG8Q8cJp2OzzeJjdpFi8RDEOGRJ7kx/bW/XfaSiXbFIgg9q4UCxctodL0yThevg+pQ9yuYdWEP5
esMWSedEyn6mbi6ylJFl9AdOLj3XTeRStRx/KGS3s/FYJYgKc4JLZR8ONJUa5McF7XwBc7dXQn7k
CN2S7OzGzpK24gbwsQamz+kG1aKq7Z+b6noBQP9sVf5/OClKKasM7tfSwAn1XKFDXOR6j8pBz+iP
N3mjF14EM7/bvp8JMGOOH8vox66C1vvBxhLkOuUIdwCcWWDGH1qgYlEg1ynK0iO02BNIwtfZBpI0
UZdvdO7HSewUHsoX2ESCfdLhNrhQqm6+onBGUp7O1f4kBLh4tkmY5Jtp13lz0iKvpz8na51p/HSP
PFoTmZzSNRe9+nokm4rMfztWjmpTcFTg6GEVDwcVT0uc9KcYs6d4LgxFz045aDSwf8Vb0yWSVG9o
WWnCpKMACK8VioKTGW3d01j+W+FBMf7eGyuLJ+a9TBDVWAmEpohtLTewoPIAUqrEmg+qnzXoofJI
VRscH2axkGR1BcppcnAdqF2UQi9SifvbJIRfeoqKQsiDaTStHm21C2pFPMsBIf6jiq4G/jqoVsyt
Vkl5tO6p9W7X8dxZvH5X9Xvd0oXg2Q2W+l94hKHBe5EvfLZuzNKEKkWadtynnkDx4O+d6K6htzS8
L7X2Z8S/leJ9u+2lPfjUyytiCEiJhzkH1Sv7qLEp7Bl+5C5bhGOyaoCzcxdzJwRuHmhJ0AT/+Y5C
4/S/aWAhbzsK3rW9las8nbVhXcRRGXC3ImEUQI2HdD8t7gWMrJCY4Wcp4JF6yCeP8M80i0nhLpj9
XhjButnl84ge2CKd2azKiUzRwcdnzybY60E2wECeq707kQWmTS0gcfxIyxKFNyYf/sSF3r9YYtEB
jU2MM5Ryudx1EjcMkPaPOgQBypOVhTGDXnzbERqhtS/7EGq6k2J0JkU+PjD0edOSkjJrjYr+t+t+
Tlv/DcWPh1X3nkV8xJb+EdHqpN9vsDVqGI4bjxIDQuLJBNoEBPfY23ehnsVYJZ4DkXcwngJNCBiJ
sTv6itLEWQPEpizGm5/28/5CGBaihZ4tMOkNW3K7AOgqEodpOeVLvqEi0D/28sI33nDIaJU9004x
HZIZOGuzugtNQMLI8tp7jsx3qZZOcd3JlM8hAP7zBombPf4VQzdWwqkBHMQsNB0QRUtaFeNvUmwJ
cfxUC9lq3auUBCnbvyibIyOQRnvCBR1p31SzQDsb60q0pGu+IG8HCiaYErbKm3fN7nVqCSGtB02X
xRDU2k5bDWBddMA3QfY1M2fHac21YCKLNkC6k6JDPYhdIGd2m9v5yUHtMVyIqzpcUOndoMVf1Meg
zV6gK1ZFO+iHTM6BXoEkMm0kVLiMFgBhOBfUUnnxXRtrhEixda3FY2ORU7kUtpE5z0veK0WNH1S0
At+TnqMb3Wr70WMwIsVULJQtIUkuXOmRqAcsFqyQpUQP0tt0jWaN2oGOm3uYfiHS3w98ygG4mt89
ZxfHN/yCdnRIr0qHRVyMuPgi1G+/9wa/Jr+ROJ5C8qyZQfkwarOBuLpiYkotgM1aVieb/7/lcL6Z
017AtGavMXnYOzH4Sz8DZvyWmUIS+CvrziCqCbpTUHpi5xkkdFAs0t3BKsj1CxDV7Sxb5NZFALVq
WmtKj4yDAnzSpJZzMQlY0kdJKzJDhUugx+v+cfGXFguRTHpI1NC3txO4OWMnAl4cbMXPPtxQ7W9R
xt6Lr9dNW04NxR00ru+BiUcu1+mFeqKH1RrBoUmWfhNSCAehiFSMBx2LkRFtJ41S6qkGy5Q6K7A6
UtQmasb8O/1OWKwxe0/DY9Vt892XgbaWmJUrHON/XLRl6SLSWFwF3STJOW0r+K1zFVwnA1qVbm5D
R/Ty/Ou00NKTquvXYO6xO2oQ3SCuI90X7e3Pc7Z82njrcMKcsGh2hs2RXehP0JalSyBCnwSlhSzl
iWqV4YQer1pMiuG8Ms5LYMCKUF9CJqwF6YUokSSOsBidGTHtPVcbAZ758FXMUE7bd1sIZ0XB7j/d
HautnY90td5ZxysOnVvP2JmFltFiC0XkGTSTOOIyMuHIUgoFaWJ4zZXeu61HGb8gZEFTvsm9HqFz
rGKJ/bnQVOZhaYeUaM6uwk/tTM2dd00g7WV8++kn1auGlmfd4BeBEiaVRBYIbpNEf/KdxOrRaR00
09wo3VhkFWfS+jM4VCsGAVmZjL987nRgMYLA6kNjY1HBhPIsYZ3KQdChNjZazcnDYQp4RvuoME2i
eF7I8/LVcuxMOv1hG2yakqjgQVhsxy9Kj0e0pVV0FRzBT+fRycT3mqsNHty9H4dlxpcBaPza6uf/
qKgS5DnsOixxk9Ls7rIu+vnUjR/fZXryb0dx0IldanZ+TVDTgM+HfhjAtoQhKUThfZS+2PcPigFH
3Ct1RPVym/FBUQASLXeg9yS/U8DDVglvnF4WuEyrJrSPoiB1WGafdXN13GtFNUim+7sYoBZZZl9l
QL04y5h60UxSlC/ZxTHnOEsVPTn0tFOwBxiXcbw1v3InXLhkGSKUc7X5YEmz2i9d0St3w5OcHQ4v
ZJaDU1Bu+VOvOC4lxDqQMFcS8RxPbunXQqF6IeGIajxmu+i6OMsO13dLN6Nijcu3Xd3fGuaZr8xz
cMTgsd9ud3og6Tg5a0puV31j/QFwoJQ7+sZ6ZH4eanJenJ9dx88ytQ3iLZMPPELfzPnwr2iudNLu
n7YY/QVIttxhsKtvznG1sqEeNGPcb6RQ/tQ8zv93JtW2M3KfGASn4+5v3TReltZvG9Mxh/gQwQH2
hJZUZne9uJu6rSSj25FslwIe9nixhklA1SYDvc22qteaSmMQ3rPqy+SHDS/FvRq/dDl7X5Rr5G6/
N7AXVMW29rJsWRRbJHpWIp67NPX8mWyVzNXrk3Hn9VmyYe743SpHhHkO3+0B2SyEwYoV24FyfTEy
0qjGGm6nx8WhMHdzAwAbcAv1NvdzNrWWxflG3DUqFkSoDzNDNifRYRJmfasFYmk0PNGAeRThJ/fj
ZNWJHgD7K5P+zFXRadtegyy+5x1mNcx1l/Hkfv4xFVUm83ZRVYEFpSlsT//XWBzSoNZe9E9IfjTG
EQr0pxNS02b1myaevFA/xTgD6fDqW7FVwfgVwdywuAJRggVwosF4sRkKpUuDIz/CGsnK95hsymHK
DYCOPvDEO/ZktTPSG0SWtg7pQahbbKK0q2wNJouYVBCH/ZhqWOWRcRmd/UsHCOAjE6jn9lmMba3f
m6iQN8fFwFdxmj8u+ELpIe5luTpqTQwlHMRBYsLDXC6GWopk4Y+ZjvqngNyVDYhy0FwxVcQ1hs1d
Iqn9LdfF7Nuax22n+3qlcmuc7kId5le0TSkSZZ1cW+ymrG1C5zJYwEhABa7gECjFvkehY2doHfYF
yDu2eR20SBrI+Su2EatOvLU+AffkWTPBNUPeyCcNzCXAiq9dATb6BE3hBkkDcK5Fxtc1G9UUxIj9
f/ZTBgDuxu6CSur56F2qrsU3yP79t5KIia+AAXueny1P4OgMkhAd6WWjlwy4H43JukrcqLwSwAeA
78EhGsMTfgg4hVjRyH+1Bv4dv6Pr31LNGhDBZZEJFRoYh+6qpDm4+avnpsge+93O2zFkkYMllSRc
u+v+De2hUESjb7pzxNT78lc1xZ4e/IQzXb37jyX72NWCKy9csKKLmVtSzTlhTwHlkwARqbYXzYif
xku8EzF8xKOnPukXpjPSasjEAuUAhuNcJRNZWWZjrO3c6MZU7YckhBW04glehLu7kuRwTblzvJU/
s+C528dzOsesrDmeK+vEOduOo1p/CCjDYqlvqqlal/InOw07uHef79miTiHLHY8/I9GJIpkHhaAg
6RrXKG0kWLaQoo3WtLKkAI9Ug0f3uHU0FlsFXdFT+AywtSW0xMwCJbSqNc09HoW+IPF2J1Vm8AkG
Y97SiOMW6ULW5gweMPR/50UzMMDPF25t/KdNDEj8O/anczYXg1r4/GtexbhIQo2Q6g2ZkvehFZe8
VjYm6MFAGMkWNabIO8Mzhjbx3TeaND/zciaFJdf3n90QXyDTL1o+6ECAjFrZrO/87lObrqbTIVtQ
FtmqDTBlbYcVTNobw+1YULLfR2o2KEPjVoJ8CM5bBIBhYWRB3aWNc1DZjab7hdzFcSs5k3X9mXDm
Xiccezg8QoVn41J9jfAV8X9HiuiAXpqqUGSrs64tlbczbhcfW4Tdml60C+1gDF6QRagfR0nVLmQg
/NbBpCpNS/enUcFO2USUcLWzdFL9p4b0Or7JCRyoCsF51aKNCFL6hISfN74skp9jsRdsBhD6UQMc
f9zJb3GTvMAJGAuPvll9s6xet7+T4wHVD0r5vd2pfL/QVUtLq5uTrxo1vZd8OB/T4ZV/n4oa1eeT
3qmg/qr/ITGQniH+Fn+GBlNqEj/6KhK3ane4AKAPoOlp/K3ElUTGrHip5vT8ZGChcWQHursWcaFS
WH6dI9pBGEuCOSHYC4TwNeQf9DeuV3i8MBV8N3ePpYyZhTrEj29yMcDC+lTMgcfNd0jz6Sclb/gV
qvLYERHY5999/KiU1kffUlHdh3ib9VIvrfKJhIZqi1yv//0ywLidFiRVjdR2TqYM4ZMKAZc4i96j
V21NqlrX1tr/CvASX7C7MNT1E2j2MnchddwsIAYpWyTM/ijVM6P+2RJzIhY3SqUDiGqZna4elh7x
zJQtSVatEOa/tgLCM24hYbr4vY2C6nSvk4gYBvC5fcovEneabOCEWRCRfppR08LeyQ/4V8GbPGnT
c7XRLUa1EQKwuuvxatSEKfgCTaePUWYrUBhlNmVAV9YdPwVKCi1yLCrHfBF8FxFTp67qWPJJcQVg
e+pjHLj34dh0MNjjXJoLViCudWKbDs9QJvIHDMvTymvbk8z91/Gb0Ks7dtIEPuqRglGU8gHRPKWa
Qi7jfN2MgFonXBDTW/wbVXUYUfczSmLE2GW6i5LjuIbh2d1jKtQItp7eFkJZVnJ5XnY82IbyBgyP
vUHf+VYaH+mt4HaIreQ2Y7+5/M7njrnTCG3ZP3Dyj7unpOHEQ6KbdSwCe1W/UvUhsqaA0z7VaxB9
gzfvD81GauiUGV8tAlaZru7Ppx4oy2QTjWs9KdTjCdRgm8W9uAekAE+mNNt5c7g7f96qNlv2W7Ip
CYg7VdyXAiDYLoHdR5rc3yIkydwdjHq09uwfTRa/TtweE3tnUgxam2AITYxg24y16OwoNWqMIK80
D+dEKzWG2cCscrunqLBjgkcaiAwinTsCl96okTWHof/DABiHOCPOe088JrBf1TpZJdgcrSz6Aosk
68wV08YKIIQBWz2RJXNNSEdlAnp/yaR4sdbcEVTVcGd8UL8lNIUsUQo6wo0h4/+RAueHOhaIifpF
NQX7maVZRrgb2P8D9ikCgPr27Hwkhe0X10uhlArhUPMcc3D9treFSYgft+VRKkQ9BMaf+IDETNfN
srRyv3Rl7Di+cGzfDZLJ8yP75rkL1nSeLKJYKyliYWCjIlunVK7aCAVFrrsX8U/KCBVFMWyO8mxD
TDiWEX3PJ01LGK+y2DgOz8WZa6u2eD6h6pvEIs2rRAcxW+thNdfSDRCgRQjtCldtucS6x3RNaF+p
RUp6Zl30wMOqPC3SGCSjz9bWxY376B+Xe3lqm2BV4+n8PZnNHRytpC9vHmH85B7s1SI1Y97VKFGT
+lbo+hNa7Yugp9Z9xt8M+OUy+HjFOqM+vm3xyqh+TW7GMhKsmTP2Ee82RYkvInfIaOmjbbxXMg3x
fZ2gcKn5u9QW1msw9cLwrDY9xV7K1dqez9LVPYYeXRm7ZQU2ihlnbfVcJA1sDMIXaPerbTDatU3x
0Dtd2cz0kKYb+woZ9PQ0MVbL2FHYFEn+g6cH7IeHlqi8t3bjKl7XQ/ePHeu+iTB+5xgmF8r/miL3
EjUg2+P1boslW4LO9ZHB3dlbjznU+hp+yqvn8Wy3/DPJF1uWCUAu+INUXn2lc85uT+RcMZNA7STE
Lofr8seGP6lOkzMskF6S81XyIzSIv+17DaruXvT2hv2H2P5LTwgFXe3qNwXienJH0az27NtPma9w
0icq60X6PGfCDA+9xL+3grtPev389FM068BvWV/jRuHPKpfQ2OQuCiIXXTmLnStW+5oUNBQcPr3L
Re9rI8j2icEtzgxqW3gLEpaPtcMVQuUYI595K6tzVypbWHACYd6XEQHzn4VXjXOKUVHHraWS3GGf
YxntZUnteKjnNd7IydAxJdnTX6XnM41rUyAOc3GL2PKOHYimCrND0Ni+jbaM6AAE/dH33QpVQWwr
klgIiLdlnba7eWALggfWm3ToqrGq5n+bwyD4yn7angHBz4ZZ7H8VZJCdcI20GECTM+adHbN6EbG/
+uodIRFVHOojcpgluxRTOXdaber2xuoScb4vDhFIGopLlqR+U62bQB1KTDMg/UdkS3HDDq//fTa9
Uoyi1R5g6yAhD3B6C7DvrXZHVylKbUS7tS4a8NuRbe75ptLmxQTZ2wzmrfP9QJLiiVYrxRON80CH
2xQtNHqLF+w3+cxAuTs5EsvOXCdMhEf4bK3wA8EBgcQ40NWwW2JrbuZqO+lpmmeWRXvQbCXcxBc7
Ue+obaClm5QvGfVFrJGNR4GQkGzdC68fwBoCaHnVec3k4ov8TXJtKeli5B7dHK1KKIfIfwRGyEES
CoP0dVIBfAMSq5TdOTsTVAEC0pqzz1VQiFy9zuTwr0FqLYnwtU4ygQGSglGvz4CmGqmKHATQe0S3
4cL03BPMgBZmj/MKGtLc0KnIpjybgfuFFp+sSABhF3T3X5wt4fI6c3qRLPQ8DbMYqzBmjs+j7Gdd
jQPsolYlT3mFBKXa2M8xsmouqzm3Ch52oDmSsuXngTHQ3sBVeV8b1bRxgTNQ4vZh22XzkDB0nnqv
ivQgmsrxH4aQB5XVrihFpKxjltWnFOyy5zLp9v3DDHlW709CwtHjIJXDSohagNEEAGvU7L9ABOXM
nnX/zmrr6uyY3MoixDjJTGTVJ36hKloz2wc10v89Tr3R7/1d6bYdVXkP6WbiQzG9W3McvRl0MLxY
I+54ZNUZL0zpwLpkb/d4kDhbLJi8w/+JEKq4gmHqu2ZNQHO04AMJIj5KZz+uUL1tuj5QzAzoGdXS
AIVVvy3b+lzipWdf2v/uavip1ciwpo3TmdpxAi7BlOIPFx0uEMjHvqG7vDFCst1qFIlbkUCH2U1g
6jXcT3JpDpuSD4BdrIEg8Gmq/p4daELTS0B/keyYt10ievJ+nyzi0DKLw1sPCF8tz9y0cmKOsDSC
VCasUlAZD7CoDLh/2swJybYYtnlUgQqZpWvST+poqQ/ytWYGfcBmWVQqHK+jEWr6cQo7d7FMMhfY
1+1zctlqwsjqEgR4KOSTqW4a0JHeLPT3cyQJ8gz8/19unCIg3xCAu8h+ZMK4cLf+EGmN/g6iEriA
Xg5rz3+Ya6BvwjObKDwOkYQ1A1c/LKxc9WHDUHbpOSyuSt2tNzNta3eXDpaZls8Pr6q8RpYFl0Dd
Sp9QnXK8Tp6DM7OqrQcq5OxIw/6Erw1ajkKBiSvsKRrPZGzM++wb7KhJF1KAenf1SeKqEsyDfX71
dmKerLg9+kdeFl3HCnVzYa0leDJ2HsMpF/IZNhmWJX6SXje0S6cPPU+VWrjHLDgssN9LNS0Emlgl
UP/B0QblTF6AiAH7kvJnZsA57RXWzCXU45noxz6BWvrL4JLlLnNnLYDl7BZS5lfnpqBehG0aPXRE
jyL2AKuqiCdR2yppMHsTZoY0sh8OxIYp6V8q/3kQirimkoFjICRXFeVC5p9tm7gIy7VpBm3MfbyF
FBLjjWU2pp4ReeK4MYcgQHGxOs2jpAMobyYpLgZfJyTNq3MGj/ZSb65exC1CYVLix28f8nElAcpc
yVXfZ1s5W8aom2uqgTSW/Z+C63uMGH1ZCcdEi0a8JkUolUtxwM6ZBqxt+I7pnTOOwP+KgZv31EP0
qaVzAk7DZSUdvg/NPr7MlxHzxq/AUk758eDjGPry7OS5Ptyud0Rh20KbXhZ7k/kFZvExxvY064Gi
TeNc2Jl1Y/bcCb0Uh4BBdgfHq8QE5rPK2VmurV1gJDI2YNXSgEr4jimS9WiFGBXR4Z80CHpjgOc7
fyZV28/jYkFOEnaVHZcBzJNNXg+k3wyzWgNmC1RR0qiwej0gF4A3GocumPV63StpKLxVWAb7Zh2q
eVs193fJWk2m9S6HHZA7I6fMr85SMzsAXOGjJZCR5qmpCdLro4SCTib8NgyqB/QbpxJp8q1MWD/E
WUwidwOywPgSOAZCcJo7ngXQuiB1TY4PWX3n9oRZQ9ZiMrANrtfCZT7samG0AchjqBV99qbwNr1J
kXuNf0uBj2nIhj763jTK/x8fb1rqqek3+PgOtT51/Ko0dAOISyOW9dhWVTbG0GfbMQoF16IpBf6F
MI4r0pyIzoHiQf0I9TXdbNd3YhtNGwaP1whlKjGr+772O/8OfXMVcasE5rLs1LOZHBlgdeCGdtMI
mbbotNmlLrU15P4Qhk2ui0DPyiQgAIID0+0qgP6au6yP+Tt7UT8eF5omfEM7BFawi6SoWF9eSOb7
qWdwdDNJ3g4hQUeHB5dYfnekQ2NQvHYKcpJPoJY8ltddGxPJGlqKsN9F/xfBjDEXjs6ZaXayYozk
t9z+kRccDILqORJ/7gbbVtpwI/Q8xqvujanFs+pWa6/6zW9nkvZ+2+NoQsGOJbiYVgPjvUU/Ptxr
mSU69wP74Ce0hdOUtuKO67AqlgsgEfrD2f9AO/6A91xEW35MNp9vSqJezmIzeCLCy/V4Aw/EebOZ
IPEUjRQShjiH4cWKETw3qbR50ENX9sZbD5vf2vtnwArQdRQoYrGFGECQHL9WW7wr1AAs9Wrp5YbE
j+EMvXvxy5wTggy6xGfgFa1ckew0vk3PV4OxepPLMzD05DFHHVhuKpX/vOpC8KbA+8qyfDMsUASt
odeYkxu3gY905torA1T4FVcGfKVe+V+pKuAOCxj/goaDgnTeOlekcIwUAUOPbEA+UC7loGK4ne1c
OzDo6wnFKuvMmm/WDnZjgO7fQ7sTg0JM1XPoNsOQt0z38pVQewd5wUSXucxlg/WnFvgY+sq2sLDO
ZiRKrMRT4BqWSKgxpk/EMviJc/eraJnY4iZsrLAXH3Q5KkzJ4YRw2Zw4CYGDC7qOqeZfW6+hcucM
62RBEi3YewCOfvHk1o2zDoHjRkSJPdxjLKCe+waqDlVSGNSO/JsMCvPtLVQ5xDvineoda+48PVOT
ZhnNAECwT8mYZdziWrpEZoYXxtoD+tzfUjCySFpEHbstNg80yc1wPMkrAT6h24kUVWCtMIKX+sHu
6og1M21Drg8fB272BJkVXd4J0lbhYFupcqeTPksKTIBRJ2oN3lSe1na5dawk+MLwu0h4FKXRJfHc
7zkm85KGxjVJl5hXhU0E2srGsjcDRGiPNWiAaBlt8h3aZuj4GzwMoYcbT6MPFeawt3MnRUtZyi6v
gJKkgryj7uPVyBjSz88d+sdwruEDOx5HwyFjyQcf2HGAzO/mMvpX35INswSTMPJJ3Gvkk3tL6rUK
SqcrI5Hb1S7tglfC/sGtE5gDi6pg7x9vibb90GjDFtLb6PstVM/wCDun9e/4bCICNw1xib9yfUT6
r84Zun7jKv8NT0jjND761tPcwRVfie7noieVTuhGaztmAVDNW922WqojR0qvhxtGSDKpLGbl87sq
eQkBpoiUtah7XBMxHHmiOwgJo2lgIfV8zXSWPep3pF0XVgpDDnGuW9WPTbc16Vu9Yocz3H9Hs86U
SNgIm3+NXr2ysRNwoaGGfWRJh9ue1fFxOXYDkVLzuKHaKMW2TBg+MPZxEj/IJHHkL8r6zoO5+Y2w
HKX5WBCtnInJBLLFU17CdOs5AJbvD6/B77OIHPEDKLhTJYsEThTkSznnkBdxCMwKn+UTgI00X7Ou
eVxj9ChMb6OCF/I1qS0+0V1eVpWSV+EqisNEF8i5G2oySH+8y4qi5UFJq20ArCeUF3/Occd3ak7K
0DFILGOab197p5+2Rbvom54LWKqAR3i0FC0xH6htLA9PXATKiVLn6bpuNkhvqcwzHR+Ilts2rBTD
gjwkcN7AEF0nVOK3H4tNIPn1dMakiJm3qSon+zBOZ/Z8+Cs0jvE3uD5cbTduZwZPk62t/6jERkTU
lHXYSF4zWto2oL+Zn7sgjroHugA8k4Vh6R2Q6fyF/4qoHCOdUczMunr8FggyD5Us11+McStn0rrf
fWmt+DZD/KpBjTfpyZmRbRu1/rwDSTY33FjPB2rbhBCArzxpT0V/cva9suvfE+GqjGl0hcdZogH8
bujVF8gbpJzM4+2VH1X9u+Hm27o/Kb7Xk69Dz9zb44JIml2WJb7WCtoa5Rnm4q/swIrkJK13580V
WHfMlV6co1UZN7fDVEVhgdJ0sL5BY9qdLNYP+WyfYnShlZxIId8HTHllpOKwutmV9NpGfQZxu120
jGLf8FifHoJ5ZMG2MWEDsb6DMcv5BTXDTXyRuUvB8jVx8DA1TWQy4uRZ8fj8Q2H8+zhXzvMXhGS1
uxd18L6B4lbFeRBM9u4j8OHOIQsw1+55Ywxt5nHAGEsiStlVSHdi7f6jWs6J5uiL/GR1Dx08tcCq
szDqOB28QRHQgZz+3Qocv0JA7PAEV0BKDAY1Vdxg0/Cwr2yrYUD522jkO0/90ibFB40lwPFgPhbH
jp3+g/H1NvcYbdkMX98WR8WEl389OH/Xv4dvuHyEb3HdxlzJMwyxpCPUHuRwfVYNotol1uxEVjL7
tb8U1t0vX2632OGxvrE4G2e0hWvyYSEAuMiU1d5Cq70eTa+7Udl2CSefRnA6LsVITrmTigM8ati/
lnM9Mg3MvMwkyLdF2/+j5AvHxI0oP4f7YzEzixw0NuUzsIsxKSTME1Xpont63G9fAv6x7oGBS/V6
6EYBgCQXK8RuHsieRtIe03wmxz5G8tUXe8MNTBvlIofV9eigzGlhbKmzqHfCS8exu7JcTu/cr9TI
NT0r2bb1Xo/MxBLvKIA/voJT0r7i5n3mW/ggfAxNgxZQoo509SFZqarfzM/6Yvck2ktZo/5/OY1q
yvakxkqTENp27H04Xz+jP0unwbfHCNVjy/qGFG90+Te9BwXdfRpYApPtEvA/KoJ4+a+Gc6XJroj0
ZW4UdiQvw4L7X061ycwg0XM/WH15yC8SyzjAmYmZ9NioVoAImzfTA0mD+fGr8sBG6fkV89lB5UI+
b7qMw6G23iJgKcHwEL0/98VkhkzESpH7jx7RhAdtQVyojE3s4XjMlHc5j9+I6zj2f1RBJqW1e9qv
LivosuzzwqTjGlWRdYi/A9TMdxoU0wzyXsnpOlIV+AKP/bkM0+FpZ6X8fMtXc/GoUafhyFFIqQvg
q0a1iCxVmNp7Uv+2uL1dIwtKNTak9fjbZAgimvKgxhhkQGK2bByN4jJbydVX+qtFPKuve1RdNWn2
Rkae2evIZTNOPKmSisZ6MDet5YlXJJD+udxYo3p6bsV4TTn7Aa72vZuZKHh3oem96E/BhAOO9RnZ
CWGXAab0+0xLFlbsi91pd1KE+ourlmQrWHU/tQDXrk1eGsm52IvQ913G0x2hQvkXXKntTGpjuWYK
RYD7HVSVfoSIcYkhxVPyGYR5948xvMVwK1Lz6/VSP0kDgAe70tV2lmDVbeega+e5rtYunad2Q/f2
6hzm7Os6/1a8ry5Qc+S1d4LLhVu18lFTJgliYtqwsy/2VftLfUwzerUlHYhDoPDqpZZ5BLAQsiS/
iO3J0DpFppdFXQA8wfBWgSlG5Zl4yVopTdsdJbQvI+bTqzZGodZR1cm+1hTfmQcZxDBJqvU6WE9W
7VLUHFp2qIARHuzll34ExGT98WUjqISx6YAF5S3jNZ5FyWoztLdULOalUjp4JYf0GgUP+xePHYgs
pFo8wHOFUGbxuLJFJ4zJVC+KWuDmNEejzextCVz+aGXkPlM9kZQQEA1g38TJb0uxYNbWruYyByM9
OFulrp+c+4HGwzCEPp4M1BVuKH2jfirxKg8d/NsXfCU0tyO/2D4Vu3p6TY2kC1pmZu9b59aRaTB8
/qL0vsMSR5Si4XYraZfvbaOw/iQCM+fXX9u7Gp9QfI4MpLrbdYWV9aQ6t8aXE0xqmZzwZlJtOXk3
kFhq9/gsNY+RlH6B2M0fdMqF9g/enZnJ50uzkFSFoVjCiiIYmKKXZiUBR6aEcwaXcAcZpxyKcLIb
tevvuPP6Q5rlBG4sBfxVG0lm8nWz2R+RziuEN+svtv6fY8wUEe2XFaeV7qyU3tFOViFwAQ7/tq4g
kU+7twrrS2/r3q7Ew92kDJHQ0rzrWQ7vmtbUfGl4YDfIJyCWqgr+QAdsmc5PikcS9lod7CQduvSJ
e8ESMpAOCGOERJPQ4yPE6QWzLM++7ZLZsGDoj0IYoY0FftmXdL1SP0gA3hCVT/oEOEfXcRRsR1ci
8RT8WtQxUkc8QUfBdydXAguiOMkJZIUWW5xCw8eq0AIsrEZY9cEjm+wNqbDvoi2evJi9A9Rl18Ii
GDUU8QlWLlCDpJ5/EDttod3PHxYI0kmtaeQ/un2gYxzk1ug7sYcyvkZkeoFS1sbPsUeZNRcJFCLx
iNqnyoAOxeilV2FBtp/ltkZmtFD0zFwfABT4DDvp5gU2Y5kdjX8RkriilaChYTsAGohsCBaxE//f
ssd5VojoWtwX8F8wkirhyU4oRk08FIc+0vLOxcf75kirABw3Vq3cRfEPsAvzslTq4gtf9yuTFshP
kFHdSJ4XQNjiW588Sz5tkpvTzppC/3jUKgtPXIOffjtusWM7twcFmW7wgWfj6Oy92jbMjHqY5TlR
HQ/UUgwZ2dd2wQONAoUHMu1sBgTYWNqdoXsrSccX82qcGghXdqYZMBlsjCe6OCU1jjm660cg5gQf
9QpivFRMRJ/rsUS/UjXOoFJHFskM6rJ05gG7iKXrjOVa8caVcrQLhjxzFuR7kJjyvD+7JF0CP+mO
nEs5m0hfUrwPXtrpfDMog21X//MfGaVrM4qYaeDaqbPOaOnosqy1RkDAyqaUPddMv12cD+EGCbif
xJ8VYUQNTEnSFwgJh1s6WcDYFYmFb4tqWp2c/p9dH7sVIXM4Ne3KxPzIdfjrHPV5+UFh/8ZAvn0r
0WeDnarVXIV/vCUSrdDLvCrR+HxRLUe+rIA46Za/XJST+oUXlHq96DUwffzZiNCuXemU4WkM1Lsl
U+gnsBI6utVFOdvRirvslSnhti/SUsH5BbbI1Vg/wPFxT0zDzmp6KK5D2JhorOe4aJiVWubFH/H2
vkUGvMx+KaWncHU4/hSwo9/5nbvjbyajRSITxKhLihQ2Dh2yZdQ6RdzLxq1awmI16BeMTJmKYDOP
WGtQttCDDUNnE7p2m5snttR1qvrjzR4WpLmAjuRH5Ateub2OB3VSQ9i/7xj6Cf7mmtovP8bTtm/N
89hRZEUsg9QMSSU652KKhqfDgOHUrYggTG2IPdreqBVSZyN4GmEYqyaPEHiKs/N58V8FePkB6i5b
qae1uetGpPsMvkQkqnP5KeI+lw4aq4evfHhI+apLeM+j2d6vz7LqjYDzIqC5hSpuqvZIc6F52PNF
PYcOaq4dDWDn4XML0nD4s3j4vNN+w1cLDQSUVEcwDwBwH7ehvpiGA3g7zhOkjb63HN4MpjVQUaP8
4/parGwRQ2G1sX2uJNXAau8BLJ98UCWWovG1GT7xv/k8a7nomMwCiyNcUe3hy2t2rw58EaLA69yU
wyO2o46g1YuArwnHzqc5X9HhR1rWU25B/SSx0LavJBj2HD4Sv3R4HIMwAFGBOrar5PlMUwT0x8OC
wvz5ekVHrz6jT+/IMAspSPUtqnd25rqJ1jEOJsDwW5KXmZ9uWHUFCfOROeIvCgErsS3D9f2w+lM0
CJ5ZKriMM8QIZnRKPmmNszKkVhrO4oFRrDuiP9TXtK+z2yNIDlxA8LJfWrd0nvYJXahA70znLI4V
hjnowuK5H1faXBaJPCn3cpL3lu+kSWcxchi7lWGiPj/an0xPG2j+Wzq/iQZY5AClz83MFL6BFHpZ
tP9Lqz5tec34H8c2Ij0AW8VLNSwmxZ9N3VIer5ec59ILyncRT/i0ba1dBz4MBaXNgNZ/4cluQB3Q
WSESLkA4FDcsypt7DLLzn2RkXK07VpG1rE9uB4NpootFyoMa+qgV6igfjSuNxK4ZkqX/zYc/ypap
OFdFpBqk+cWLDZ9jAL8o8J29/gzaiiPEmv7ujJY7jhUaSBESrR509c7xjjc4mC/IgBVlntfNYJkQ
Mf8uTiTNI/SbzK41C3N2nTwdg7UC6HYRe7eJa3TJs4410MH6XuLenczIhj+fhcvH5n/iq221tp/l
FIAEMDSKiAa/Ga6rCusQrxXADzAXbVs2woUTHDFlQDOzT3nvSMChijMkYGGDxWg1stUDstaRUFWw
GWUdkaKgchimcB4MVbSpLiEJCSOaZygzBX+fHCwYDm0t8BDHEIAmb73IBbeBytcxa01qUr3EdkAU
B6SkyroshxGHfhwAJf9WW2HX6OcuON7GvYWVR1REwwo2Cvx0tpyhxIbCt8bwffo+E1Wkq6LzWeGd
Sg7qw58DAcbqXBoZD0yX8gUvVQJBV4L/AjdPVx2FbFdEAf2grQSbGtLIy2WX8+ncL3YdvtJ8/VjD
bXJNQPEAU+cdN833PZkOx2w4fzys+UZk9LeixHneJIQ+SXTbRt7rHfOHkSOsGMmenJXadYtprCiL
lg17nNlnedHNPpYR5xe8x661xBK3SBx1tpLisacwOu7j7MBJJMBaKxrHtxUr28/2K7MuIm/h9JLo
7acTg+G+S/wvgqZvZelw7nzRGiSxljn6n3ygU/4AZxWOpBQe5ydPoNcOpefd9S6/IUfL3pEK+okx
pMYjMR69JluHjfO79tYo0mdcXrH6XFpvY6EUCyJLHfAe89Yg7hKvKnV8vkgHA/Wwc6cRooC/a4O1
obw6mK94/WJiLSXEBRB8MhE5mJnvjNsE9PROVebhJITnKJXPHUXUrQLjrBJFK5dDpyReBoiekIFT
gYSLk3arrZKeYbSdgz+ZKIoZw5bSJtuZbadTbfBFH/eLjhtRNUlr6JWf1c8EHsnxbaHQ8C5mwZGc
xOuUQpUiIvrkIZVrjJ55RkLtdZaVSFvN+gERUCOcmtqB3eL6MEiDkPvQNNpJIo0UqFwW8gegHKsw
2u8HyWd8V1CN9XIJ7OJ0IpN+Q7YJdTdnsZ1a5DIGJbnXH+DKiEtYPt3Zv/V1a3VbUpjQSdjRmidn
obpMi5XuRDTLq2/t/2Wfys2nrOvh7weyXJ2DfKPySq+laYpOC0J+5gV2C9ICkbv6xbvrfQmFQfGS
hCjgcCqz6/QE3vjGcrJQV7Jgg5vY3wry4ibJ/TPEtBHul6k0n49/PzCobWsQXN8OZdeq890T2wDq
tF/Vk4IvFbun1uS4uD8GzFvOsW5bjJNiVDnDEz8NMtF7U79Yzl2Yu3I+xIiGxyNXVfyOo6K9eBDT
PLOOnGUNII9UL8HfaLHwG59w5xhdxj6rSLHF4tsy8et+suC1HGJSvw2DudNzcEDQbp1OF8drtF37
r1d/I9ERmT8xUDMCiNB82SshfzVRyvUwHJdoCenYZyh4ImuMunEZnUx0lCK3KjlBxVmXcOo242Ll
StooZGfYDYrI68cEYDkaG+HF5CJ/V55PhvBKT4pkiTIArnJ1Mu/+DuatupZf3mdep30XP01EeWVi
mRRGqUG+c2h83+etodGkqwwbsxX5pN8oNIFa7RcOiXynm9d3z3pGIfM+k3gPGgRkbvCg4v+53B6P
IaNv7UQ1lmgD/lgEj1sZ4a0nswPL1cazACwpQXbBBW6ogjNM+YnZDU6Y5IbNq9PKPiMD1AkeB1bn
SS2rPvCY+m7FJ0Reg9D/Dx3d5tLSlgFceGBbO7Jwrhl/dq3276BPQBKX2dmMhZXeYQHMwZ2eSvAS
ZWV7GKP9mxQsLT+574fG/0GWqjjs1EHVJtLZ4MSgUpNNPrkyXn8L++18WGRBkAS1iUWDOpp6bBkW
grYw+aCx4WnOfLVCoG7zSMvH8AfC2xJiiB5MfbXAnw7Sgh0CdkrASpnthmfimB8kAAIvr3zi4R00
x21OuQqWU2bETL6mpemWCwZ0ppJXA1UYLv6YzzZt6K1l376GvX7KOQKdM2n/bMM6ZM3N4/jNy4El
lruhBiYlM8yO/9Y7zTGhuIM9pD6u0XbzzKh8t84tj0+6BIAEcOS+w7z04XB6WieJ1j71Q6UtePKf
KnvqTX/+4my0VFXgVspmuZ9vXdgMAO1CP5TM/PfeDiTdcoR/QcnzMqe6eOEGXP55dyYe4qycgvPf
n8CMirVW+CF46Rub0LK6+mYQ5EvALX3CxWMcK1U6YgeIAOITCccv8gMnuArySZoTfvs4ncRvSK7B
Ha9pL47hRH8H8yJ7pd7LthekSuHfsDBDanpuja6tB1HjW7Zx4ur+uxrgJkDU59mEQH4VSzkGyBZ6
rjlpHmJrGCcfYv29+RlKEG3n8DIhrG2qoi52hGuSzKbrN887LLo8xwoNkuy4fWzAJypw2TQvzghP
zW4Ya1zoeuCeM8s6qC/rCwRQ5nY5Kwl2DYS9+PWVia4NO2zWoQ50eWyqk3gP13KhjOcwMlHxolNZ
1+m0yEv/XdDOjsPq7Q/hpdmI0SSAesXkVBSYMKVjMOhxZGHNgobdWZyqwCkzIqP0v6fasN+uJMFi
PNKpbCja/nxYtimwjbybrIoVKLgUPXZWmUVAAD6Bbuu4E1GdUCCQYkX6y2zNn81lIEathAEd9AC5
Y+nBjFJzgUIN3xVBYvKK8FCI4Ct9yUX84ijlbeywtKUh0oV4BduVrdhXGEcLUkCt+33dlSv0SPME
lAaAmTo19Hn8fUJslriKM9q+YvOEbjspqZCeQrc5qNwLqNW5eqYO7db6oDojLDGozT7Ypic/PNC8
gfo7hIvaOPF9Ysp2AdvCRSO2rAOJMNZuWImatJJ3uJt7ccQmSoj0M8b95Eu4d6Wvf0H4kko1NgLD
TOhmFz/JFdVAIt0PwfVQbyYWpaCGDxupCtgSTa6eqfjMpJ+tcHR8LcedQo2NSsaW/kv9acEycS7w
aQwYk7VgFDWo0B+FTpFLJd15DK5fI9YZbNi83fe6eE5Bcvi2q+JirJP24c5bXiVH/Q9WQK8l2SqV
CYoDAz6hDf1O1dWvPCh6G8jYYdeZ62jQaOTEdA0sNSWTCw+BZmUvf3OtlA0gIFmyq7i1CyPYGKOR
jGHhXYzmrEGXFkiCKjssRV1gZ4oMseP8bcT+vFXLNFVe0t0APJL9qoTeoqQ8wQnNUB+GORRpJFOg
oHybNEqIJr55P88MoPuPSmAf2R/4ga5dwv0shKoB8ctUV1O3dfgVopMpZgDg3W7Z2GBHb0NnZ0Zq
4biK1+jdJCMPxfqT4TFQ4ZpT+7M6uysQQg8/e1FNgTYycCBjy35Cq0gmJW8rwgPuq7EY3Nq7weL3
c+L2jWtyuHD0FgiJj6Wa9Dcm6KBrVivVTkiML5KONCRNtfxMnZGuPWEcordVhbt9K8knzhZep4gS
5kiZ8kwvZQpYRO2DKBde2br4AVVYYZkGA6aGS1rFqZki2G+Nl5PZGlTmlZDhYcth7Kut2jeXNi2a
MN1u7Nh7JSpRODUNnNtHQY0OnmYeo0jrM2rOOraQnQ+0AqISWRlK7wTF/PfW5uORjJNMZQOF3NKu
TO3afbskdf1LY86Hkr50yVQooimmHdldY1Dva6bKrfjybeVYcT9FPFTHIVvmUhG53Wc7XjpZ98wk
fqYMtzkcp4flfH7hRYgiMO+DgxBbMcOamqawDs/db3GOYsgZ1rLQhfAvJ84IL9FXIF8H8PnZqg1K
bjIUOAsgN+oXTaERhXJSIb1+IWnIrEftiHdO5fr/ZYDb9MBwxCKi7LMGZBhfLKnGbkOps1cH0fsx
a8YVtPdk/1+zm6rFFj0v/4pNgz9wM5wCKiNo31EPld3Qxahkyr4wy06G1NqcCM+7K7NJhTEJazst
XaPakB/WCDYHWboZ4Vnr62uFt1hwAU2VmxemEDDpx4B5DmX+Fh/cKGm7C0/MtzkbGCVvCMCOm3px
BxUEzvdatyhnBVA5olXX9LzqVZ5CFhQjkjwYYvIEJQ2to1Ht1AJ/9Ig+bYM0qxK8FmcrtPhWFUtF
WMdmYuA0APXqQBz1WksLH4scIcRa+wiyLwWhfPCub4GE7a2/MY0sXTwFPCahsjlwLoZvOg80XnQq
w81X29lF0V6QNtZdxn6QzRlsCKpOUup8R//xMQau7tM0FXlnzylhOYnquB8CfD6a+nlcgw9IrrvY
Kvxm4DHXuNG5Z8E9kWtZno0vgguoVZHQP/Yz8H3QZ8HLz5aEgM1Ryn7TpWHEK0b8OqHhyvDa34A8
dsk1/X7FteBjvnImHwSQzIB86P48883LFdgbXF7ZvxbXKpYU0zm8yYVqztG/ScI7qR+RLF8/txp6
wuvmHpzeTuJ2VIjJVEcu7w5xoHd391P/Wq446ZFKk4SoILsk2EgL/P8qO9+h41TwZMK/YV4iV9kb
ko4shaX5sGQmaVVaxsEntC7SYdYyl092Mkv977X4XMiUkisIXeOFmausoI2u98VsbetJopEBhWI8
U1cE+JFyGJMS2X4VHLCeVXQJcMQ7q+WaBw1y6qOpS0vRp0PLfeVKBI1MLg1GY49/tWks+rN0Db+x
Zh8RkApZ0Sdhy0XQZeDFrxW9FDDZAfi8rerTXxUpdrwlMk1O9P9S76dmBNYyXdwmf8Pm7EbeGTuY
oxbEg3Wh3ykbCk8vRUWKy974TiVQqyPSrJcJnqLG4e83lRHcf/jIUV8WoFlMzDAPJNvANYlwZgj/
cACBVAf4Obkj70o7XjgHl6CfoFdD5Vl758H1iFZmyQW86Ml3RidnnOK+Sa1OSrEd4zt1O0VoeuQg
oeKEGwf0fJeJ1wVTYCfOclzfuUpDBEE5weUtspkxJk4urnoMWdx9sQKoK6r4cOj/FouXM/utK6e4
oMdPCkuj+i2R1cpgagMiZaLk/JUEMhBcM2BKEcwmvhvJ/NwtTRuY3bllIvMhGeqxvhXLODrYLb1K
qvR05FMlXk/C7nSxvuIFdz5ElcTL69YivpPW1vNFrWFjkWGrVJlgpjOAGDxzt9eHbYMwGZ0h67fw
OL5AUj0lfbGaEhNA8gXZQsHZqOhkZATFYNcy+EQ97NKoag10MeH/dr45ZaQhqdoLH7cv/IiwaIqX
XSNeEhagXkWoPRTb5W7ugMmsUXKvnA4j7U0JR/x0L8o21yZNKrUlhs5PW/jYX5ZAx3H8ZvpD1iBz
+l+6WcKvxx9x9r8mltMGEGxWW7YKCVZHTgDrSrQSaj8sqYSFq1uihOY5x3WZi5mhGtMKldWgr5+/
iIfeq+3nKWe9AzTUHAmXNK6Y80QqNThg/9QK2ZhD5F+qH8ynrVKWztfsLZd85sSIw+jxYaXwMXEe
jzt/Z6i7ZnyED50lJ92HmT9VXfH8GK/PQR4J+QNUF4oddcPsfqO0pGjIodzCMl/9dxSMs1m3Udtx
TQaxcCZ/Dc0VEwEh3Sj+zZ735gFFCzOhxhmB2Dws+CWKIgqi++6lwBvExSHVAajlg7CbFmUebM2F
aAv38MJltvLSjo6s9508ad/FghnnXWStUFGL5Pa28Ul/rwO8bRoFd+Q/YDXtCvBJaPSgUc6JnE0z
JxJarPIdX8RWesOv2Nhq25AFOSkPdZYzY7MF336XkjQxBZlBGRnGr6UzAIBBmYGIwg94rJ5RyIjN
fdlTWnHkCq0IHEUUFoex3XXXQoFbMnKbdG2t42ucP6u8/VHJJfNE2NYKAJJSPzMSfhi0UfssX750
eF5RQaj8U3Q0imqzg6Bt52hK3oY4mUuqcMsbPIbGa/2+dYQBvBd/Xj+w2RUHvFm3Vx1OQLGnzk+d
0jT9/BzgkcrS/a5JFqsKOWsQH5Nx0H0QMJ0/0TQMp5lPoLit80ABI+eVUKBVCdrvMWHFb9JWoaG9
hyydYm5ZlG/Il2BIW72fPIruV8jr2ShXilMZoDiLLEoVOkp3RyKzQrpszG6bmIcMOYizIq9wxnp7
aeLDYcnWdTad4ahAxInZrWBsTQG7zZXxEcTuSlds1P+29oRZy8woVtCae4hxTWli84ZT2H8+pT4c
E1u0kdu2bQDlt7kt56fBRChNm9icf3EJ0oTndMGoH2Y76GC8jh8h4knOHj1sAhK7u0guI52HomMJ
ewLiec8SD/aWNQelYrb4RxtrP77Kno28J+J7tH/DoxSU+KfYdTs00f2Sq4cDWdYC4NMq+cG2c/2L
ER5GqP9F6575LR2nUy/kjRV8cqqoLvkjvmCzxfoEOsjd8/zIZkgOhAQeOuMbo0ZFg+q9eTevnbg+
7wJAw4lYY90galo6P6UpAymumzZJUFEBvdP/sW7+hq4jtlBb2JttKHD4GthjkJ9Bcerq9IWndpPz
7XObHo2PkwiOo05ru/mO156qmhTFRdeLwXF3bqb/b7+Rz8hiEfu/iNQvMGIaxvFZa2Dij0ERDsvN
AOMOAsklyuOKKjGa9eamtLhK3sORFBd2SMqeZVA1YV8ohg+nzsAGWdiMs1Sff7J9ETa/0pL/b157
DgFiX2cfVNStB+c0547+SgaZ/DNcEgTSM62aYdsdGKIQB8WY9tb7/hHy/MNKulgxjgEMalz98zch
nB0QYo1q1ZTrfW30OcVMAW3G0FKGC8/LJRUTeJ4d3hgfN625QA/QD0usBiD56roMIzzxiJSAbmYv
aS8U+MMQWjVO/HTaFH9uH8mfYWDKD991jnPSZsWuQ3D4SnDHItSi4F8qB7OX8IM4eUVgKXHNckJX
k56qfh20zn0ek98DciRjUUwDpfyomP11cgw1Hnol2I95oXJIK91QF4mHKy4aoKpZpwBLKbckKHa7
els1lyBH+vE4yHA/+KjJ0whtUugwUE8EWFFmBmZrZEKlUTjPw334iJ75oExewTseFkmHQxRm6P4L
/xW9FzOtpIZRyuyvfFLgZXoLHvIp4dRssVfpYxHaQstSv1Fu6s0gq9V6pdj8ln6FZywqetrrfF24
6TZRux6Pw/3eVbK3ejNe3mFQippAaNqWeG9nLHQ1ZyiyPW7mjKsa4v/J46Gvd2ILiLJ0gAv+0abY
fU3Q6vgvKUzJ1MWg34CJ4AO9YcBZVoOSd44KCl8O0TZORtQiA13oEW50tz6RmVH/MLdnUch1oiSH
Ip4R4XAgCFBo+hEbFnQQzPIFgx4AHzF/svwAaEnuILN6l74/XNx0yV+vYRkKZPAasxFrsBQX854l
n1Deb1nxVNPK+Kk4wOMNVCAZe1n5c0Ok8uQSfq+2ik7yAdfuKt2ZeJCqPksiHr9LTaBQozwYTfkE
EfI3j9Vb9ZhspCxxcSU9KwSyF4pEMByGUxFWUgaFkTm4GrMfr8A10qQtc6+Mzfln7F60edJhaIsr
7/xMqHg9HsLHNmVa8QPoHgkta+BqJHagV4CjfQyJAbGux4KuQkuDcR7xqsHG19FLnxK5bl/fI9Oc
iHeOcTi6SeB5ptBK3uC2Dma9fQ+nrZKFwldX+SeBtn+S9N3vvEgG9P6dKk6f1C4NZI5KIpMa78BW
GknxHE1WlHV5xSDBxxFHpZFsHiDpb4DdHixhulNdb3bzslM0Fn4t609ofGhI4r/gAFQ5ALMniEqd
IbYYxWr8VH9CcsMY9VM/exvaSdyzrBE/zkyOTpVchC24ycufE8RFxLCrlHh/mZymDy1bbxo4cCEX
Mqn2Y4RdzkJMceee3/9yP7MfCj15z7c4ANgUNzEVR5CDe+JFtXGv6Jxafm5HOHXVFp0J6nROLWl6
zJkXqltk4BTDaCfrGUfsFzD/vvtNTzHe1WCVL4ljPwJ7WmAIg/5IbgrFZYHuzpsDWY42mu1OcWE5
D2jMbgO8PO0bS0B6jjuWTW9j8eaXBvZqa1SlxqBUkTSvxgtdIbuFgm8YCDO3Qf+vE1MaY4MFQEmI
G7DpCRIsECh/6LBhSOHIQBW9xsbAvaWWRHwnyI3T4XPphGJN8qyXbmnNxx+Rw4LWisqlruvR9mzW
5WP3VxtuKitH0frrgIS5DbZBYsTyDXi+dBvys2UjeOglJQtK55yTE2lhazhvpYMrkmwjP5ZaZ9S0
1+U8p7mYh9m4yBqMdZWUhBhK+jo6iCnRPO7Q8olhetvngygkbffbp6MzE5nwBgu1gFIQZ1hFcoa7
yc2shi0/WYGaa5PTCZxLrj1eFehuZz1UcfVduXW3IxH0t38luaRC8NAxgGc3cBmhr2IKQo2IZpO6
QCmCgzErgs8XZAJLaRyf+l8jljV0GdMhFObyKuxyolRXuktk0VD4TmtLns9tKiC+kE6N1aoZiSS5
jMdUehUTBdG0gVOjamADym1yQUyFpNHOXQHEaPPmdTrmWrRGcPTRQCet0GxJGHdMqlOdizM9wNnL
GevloWaRDbsLvyZQxjQRMpDTbpb35RBuJS4zU8NrcmRQZHIuzaJP/KUKkMZrnuVMmb82zy5ufBfB
/uVKq/lb8LMtXM2+zYyK26YYlGZSKYONcsr4zhup+PH0TBJChFxffKhHQ0SrPaymjeTKHaeIOGUJ
ue0wTa/MmLNTXJifKZKzoFYh+NrpJJZp2Z4CjCBBFlmf04HgbszdoCv8ok3PEgaB8R7+pcYzOJeJ
ygDFxplqQCynsSDuatg4WfTBx0vvpBEAQ66da5pY6TV43Ryr3fB1nkuJ55AoJ1ivYqgO32SsBzJE
zBMnYE9acvZnsrQ5P0ICwgvDGGAzKgSo2Hxc3amXzI7h8nLoSyLWU6VGjpluSP1G9N909FByc0iB
699OlOI5WfHXlQBSnf5zPVycNP85NufAaa0K2IOXd6XdJukjXIFREfgCj64o87df41A2tz3XYu/h
XloUjl15D249Ew0MdGz8hrGB4SC64H8k55CiyeEqFhO2EUo96CPBaUcENBTekERihNY0caTeLpHo
igqBEavXh4uqLxWKwdvuHgf9q3PIjxi/dw4yGLNjRqeFNoQB79US6VMhuU1cTnl53EiPUJQvNd59
53xFrlHRZZlqIAssv9hiZahUQC0wb8esfn/oyHftl6eRJgE9m4b6qD/vFEaURyemLvXbw0hEVaC4
TczTZnYLQFt/fJSwUq1tpNP/4HOFGrEqpmds6vYcyqMcE0rIaidpEOsv02IRocap0MeKGaUUmiES
ODGGXKmeRewPs2Ng8WxWwcsu65zJDqIGYTYRAxLNYiv6vAFCpT6/ch7WZbtfMChKHjTUYL4Sj1cY
XQXTIpA8LtDNAoFi25rBGlIU0Md2RHOTzo1mg/q+2GH4IvBFA5IZWOxTLgBsGqXeVbRB3Iy+bPHQ
YGdOvlfaGFFZjPpd00wVvz1uZ7Ot9Fbd1V0Fs0u639aj12s7ESMWKAFqLTTxZZtENeVum9z7Rriv
CnYREbqQ/wAbCXHm1+KaB05UMqQ/GXrFeWYAJUJv9N1b0Y1YuaIr09YxRHmlG/BTlzva5NAYoAyw
m4kBf7AgVbkSPFnW8h0WmaE5wOBM39Eis+xDayp26KVSiyb13fN6W1+LmMb4mX6khOZKrQiFE7RS
NibcetT8eimhSM+UYUFi9g+55ed8EDjbdL+qDXQPI11gY5ZpTw3EqKSnNz9aCx7h3xVnC2r6oP84
KXK6RVcHIACsJrqJmvvvG1WpOYZEWMqo7L8jZVKXQEeLz33YmoXRmVhrl/kZk55Ab4dqZSonZeff
F0Rvg1GlKiETIbm1E4Ggxa9JA5UBH/z4A+9aJ4+OirhkJlynXGNE8DcmcDjsvTQsGVWWPZQFF+6j
nFmLu9MYTufoI778qY29KXaR5KIY86g4R8oQI4Q2RWWZzU8hOsQ2ufraI0D1SbADNirxH6nIiLQH
l5G0auLhVB4RdHrCfS0d872WvDZurVT16fCzv0eKf+k5Qz6fzXaypiRhR+1Ep95u5qARqkBOkJfM
6690rmihrzSUGw1o3u9mcVsT8PpqTBcJA+qNumcQl/0KrTCzAcgcQFFZSRYChJuhEaLxSg+3p/Z7
oXldTrWKLjwwiGAgGALaPfN25QjBh3zQuaYIpnIXIW0hf3c3iaLTcybhcO61903pyPFAC5rZBPmF
JQamg+/43UTkmN717708166jFZeb8pcXQysOZ6XNrnqgn6L5KNlxbmO6KM1s8rEqi7tCO+aMhYOL
Qa+jjP+AyObVXo8RQ36lb73ey5Ax5aVstXv/v//mYN3ayLqn67SwBSvRwV6gG/afe26MgcJYb3HB
GpBM5d2Ku20bXpkBj7R4aFr8ktLBnQ+r/GN4fqRGjdm2kzzQMgPqeBGrxFowE8AqeNce9i8il98N
hB9BMjLrkJoPCGIkJj8s48qMgGtNWYzzsAsP5scJv14HVBff4IHyNyxUfUtCdPkPk+8BfycS8YUJ
YIw9AZuAsX58tpX5i6ynFblYsHjd/mYCKVA9kp48x4uL5Gskz2G8TkPaOnnMd+I1ShubxumjUgbR
mPGP8r9LKSYEzg00jiv32fOUbStJnfUxBShaHDQsptSSOLG/OZmgNf4IJ4zhgT34mwFK6Uv26u1I
ZB5ItV5NoVVhchRM2h27OcUG01rZoBgvVvfWps4sd9lkrz3xGG30zM6KB//tyo45Ki0rkvmt8iz9
KM5uHitJe3bj7+h1DrXBWbvrigJpJwPXNIT/g/Y0dKxU3lNRTF7VM0qEtF5ndfPrt7bT/irl1YO9
T5+ayjO2NAz0SqUirKDEfDKauqOp/TAY0H18Fox92WQXMsZsNqbUCx1TNadPFpuyk9bCDiva2slo
7mAq22AWdamfdI/6e3+4LgfpBUcTGQAW1eaR7zI6hYfCYmK7TSABwt1PDBaOqz7vytI/u4L0cWBf
3hZ8K7ncOoXvfy4yd1Tkqk4np4WhIrONsAAE76q98cP3iCUGQmK24y+bzN+d95WUlMBGwrFDSJ7G
hQk2iHMeU+E1nOd4GOOLneLzYa9Z2MBB5TzX6AbFjj07LSFfhDN3Z1NnxYbGQYLO2f7/mZ+cvHxN
P40OzN63qpEwirtEWc/h5ftvkGISDIxEXlxEuSllfxKd6EG65yyM9VqZalRLrGRhjAOzOiYKVHiO
ijitANu2h92Lw18ZRLR6WXt9rj2zemrNfxlFrUXbSrUPXRn9ldX8Y1LZj1rkqsJVqRdUR1s5stIR
2uEpeI/G1y5Hos6PizLz+dH8lGLt863o7EkS03IAtwrDCbmAcSXc+Kd+PhGE1Q53V7Af1VEyb0zE
AMYVcFMcUtcVQn8bBYtOG5OmEnVUdUPGAZaOQGPqpGe9jn9YqUZ/LJZMjVn8KK52IRvJmMeEeMQH
HzsdkCYBBlHFj0ydMxvveTeLl/r345Qhptezq07TVFwDgN9xJRwNcuJrzHSvxLU+96luGZhTrsHq
lqHxg8WHLbTvsbzoqm/fDFOhvZFNmjNldw3b6MFrWhrAcX9OJebwz6afchQ675N9ctYV4YlV4QwK
lmHwgeq/+WqSl+s7YfH5VX8g+UlEavRFwmTLMsWpkaNCbxjtAnzZM4ne4sDRoiZr/KAixZrLyrY6
4bXjVtpHhzCAUvpkMtMsB9NwvgPUecpfmn9kyu1Bn8eVH38AZqNnAifO29v32RHi2eqP+7PLZd/5
irgZzek76vlvc8GrDc9X0xzRXu0GLl3DCnisdB8LjFsz/ByU9FX/cWGxrvcsWDBNniL90BaZjpOZ
JVFM4QGAvIhMYYMmht+sDWoZDW4R+yKJS64a4FQqp9uaAjOIYM8eWfsr/wF4ztuHzSPjFs7BJG/L
B9kkBKJEKy6ec3tB6ESfQv3+oqYqGdM3cQe09U2MIowMtZ8X3R7lITrbzv204XYz4VKz5v+Sccym
65ckdRI6mPsUtA7LAXm4Pvu1RZ2Fp1SnJ6i+p3hVWoTZFu6Kmi/E9c7bnPVaVUyHkz+jzmgEQROd
QViD9VSMCiHE+RuHCvsk0itph0jLTOGWv6eORE0fe1DVN+rrq0ZeIJ4vXHhnCj/23f/J1eOKz/YF
BXlxrhZjSt6lkXI/Wl4ThMdymCba2Los2l55FGFBUq0UrNbwGuj0bTJo8GdzJHrFwTDE/3DOIMGw
zT/GuZzV+3lCXtPLKHJKWo1yB795tinrg/LnLUJ56g9yzzk4zBAh2kHgeSkmTbzrzJeCo7rCOWUc
BaXk0lhI4pC8g8OxI4RNcH1xPhPf1GOuPjivNQq283/ZvX+bIIC+uWuihdGrTqOUQFHNtImQVjFx
8+sYs3ygKuwGzr8JjxOvB3h6RMsaHt6UL1bIvmCFlasL0Nrd0tBMBDDxTsifh+Yx1nx8A1jEycDY
XV9BLPJkp5gneIRIyjtw+5kYOh2s6l35XLjIiHg/Z6sCpUTlLCRGvVeC8KE9C1ScPFroKnml+gl0
fzGMmQDzuyeXosqKf7tYwrO0tSn4rFL8//Eye2S7pC9SaZ6Kz4hCml+xG61kesZU915oitQMRTdj
j1JXAtGeHIYSG+e/wXTNqYIGX10MOH4IjbOTFrFONC/cn/rqU/tSapteHeFvNBShveF0PPyG/TOX
VSjQCPHS9toyuZ1g7TQeuI6Wnjbxy/OyDY43UJe77i+v3B4WMs9gPr1nWQT6qUPVO06DGwryk3jK
L95IiKdFp3raJ1hcOuytFpSnxGAjMq73a3SqeIuWavF/SEi0r8oMik6zFM7Zn0INkHjbr4vJSVuo
ZM1wiw2Ejt4ZUYL/Q54lb1YhoNpUblae9LL/6w9l4qqi4cx2negTSuT7mPIw5G2yQeqZBbpdptHg
CTmgABCPYBYB57dscYxhOD2qRnxWA/9997wrz5+kjr5phyuPgMeZCfkfArlx03uoj4IDFExYENsU
u/dn50vqWxCL2UWG+1mf0tLEXuHKn6bL70Z5aMWAOvi2bqGJF65bBZ8i29pFaRv/OyjqtcLBsVaV
xnFAPUNyJNSd+kUpr1a3tm1eAFQZNQ6Xt0jjOtA4SMxRq4qfCq08+1NvnWeZ57S6afhwwHcsgr+K
hV+rjkJd3aH44o2KGdC5zfdDlYBIHvMQTeXIBf8+3Rk7aYHd5gH4K78xRV5utudnAgPpU9NNMm6i
RYbLWxFhWxR9tW3yEVN+YjWL2nKZP5TLfNWRcHXBrXnBeD4Z5L/0ON3Mk7xb2JMjG0BMNPG9Qg73
tGxwImv8IVXNmN0qk23vWlqmroHqJrk652ts0LI8FjRSfaQciDaKi5cq9nWhDx69rV5BKpNTtF71
zA2+kCl38qLTEj69sOBYKrEv/8jE2KoLv3qZu8aIGrmiw0ucnbZiRulbkyyWIe9JzlH7HLHVCqhK
U6oN+LGlGIssGXE8SFsrtmHl6ZGNtf5g6UEhYUmJZVmXJpvWMiR5jDe5oM+RbQ8W9vEMV+hrwh9f
zLJwhZdSV5ebvd94+VFoImqtJQ10nIUbpFDVlsppPO+W7vXCypkMbsOs/uy7qQ1BR2RzPsuu0CoF
szTxSY+gN55sXQEXfGq+9E2vEhlzZ/M4VXFkFEmJ1xY06TeGQIo/pPPQtMHYjxLwIapWeqGOFkMJ
9JiqPIknjYaShrRhr4bFwnLtWnfvFci6jwH3r9fFuQ7ksKetcwXFTStXjN3VZVzAmg4qT0S568Ao
5qHlIWlwx37OdMCDzmdfDEOnaz1ZIQ5Oq3q9hwX1JGKDAp9q455gp7mHW0XfibrZ6GQswQvRQZzu
pBo6ykuwSqMo3ZajEtD7/DDSvKTkCWz3v8q0+LKk5fT+dtj6tKiChKurJk+lJH2hjjfDs434Kjt3
IsuhHfNkrTY9CCkJF94qsfz1SlHK6t8/E06IjSvf6xft5zEg49BDgnlKNGojig4sv5D8W6emWyO/
2l6O/hKiqV522G6JxULxrCmg4+b8zK/7XNWo/MTBLaiABTZNT8ApBIR9+9q16o4ocEFhnWIcs5um
soM3mSVjilqQ4kqMcDE9/056GifDvYoVR+AOtFQVpJE2quesP8CxZVRb9wAeke4B8yl3Eo0nA16N
trIXOT7/kMC6bWQTAdPuCAuXkoV9UNCbmoAoF/ObQZpr1P8ib8SySYYw3WtIBSeVDfsgOMjvt7Ze
S2JEY+1TtZCV0g81C1NiiGyRHgP1/gULkdcN077N/+du7BtS4sZEH7PeTUVjSxh4rsmc0BpDiiD/
CBQEpUxQzBcNpTdmRNtSY0t74EmNzXODk5TScZiymCZNSJTuLBaU9rRHB/7P2+ZsQKKNioyULCKs
cjOkOCQnra20if5VBmeqjAb0rxszzk+c+A0cQorJxVsjzZuU3Tq0ovIM3V26siVHkNXLcw7ZBeaR
rqGwH1+BT86HmMNu+oauwqXg6QIx1FcbsArN8fTz2aKHlfOfvIgBBePTctO9j+QBKIIQz3bydOXM
dk9+HLvh+oRE2i9qzLYp7Md2X3XP1RlmyYz1OUYCe1bNB1/yaFfSZPUtSuu00MFiIGMapKXxQ2yD
tDqSBmInBe3p3CACygCSxmJzno0s0FivtIt7QH+E0vNfNLwYYnxOBtJLt5GUiV0aw8TtI5doLG8X
aeU4YeNZBokvkpeYa461jXxsFRkGsGRb5bjeHR/44lFcoU5ROqYcojx5NSxTt7BamOHyMABaOfWc
NyOvsu+49U48/bbZiRJMsh92nYZo3rT1yeRY5CU5z0Om7qSXMVCFwgKZUYndGLrNGXPGpELxFVTC
Q5R4PaCpWTEDGxZY8z3I8FdLKxJFZ27cdazUv3REIiL38Hq0nkDtc1PN45vDiuLpEPWWhXHK7bU2
6DZojkev/YXfc+sLmtUumu9wfQqSJW+RqFmaUMh0rmuOkUoTK0/Pwqh34VNCzSdMBrZK7GmAxEhD
CWLTudhOH2RF2AIkHHncSziv47JCvBxlfTGIjXpmjMgmAKOroUAo9RBTFPZm7vpLvPyyUcMhBBFp
kIBr1kmEc5lvYBYEaiNkUOfIDF2yl08q0uacSAZ1BNHCaHgCNTGoDxGd/LBxS1VoMDbfZan3NgM9
YhgQOV05qQYbcpN17Z7hIiaW9PInAqoC7HGXZOHfY20vygFqusIGZroHU7cbYXqqhvaphdJVcUch
JSZaYNrrbEZim/fbUvJIv6XwNcQnrRwVOc2JCwuHmSVn8JEO/1yv4Ksg1ujlrUycfX+tgSOL73Bd
wr01hN1Pbovvk4yjDFE7Z6qz3NI8NWYsh0fnie0Rb3RaHxeUMIBqGcYWapjm/Pvpuks0PsFwksc0
OpCppgVbQUfMkWQPod+eKTbG1piXEKX3aog1P2Q6X2UUQfKtDSBatJhceG0b4QFCLazlklPI2dj2
SyibpR6E/09xt0zIJ+wxvKZ3PJBrnNJR+vFQxqr9kvLS0zxOJ08tKBVLhVLGn1iHaPfpB8xCsjjx
fJ5cVWuvehYt7/PPmqjojWqJ/g4zCEDaatOYUBIPSD1Ha6ttvekT7EZgKExP9qs+kU4NLslAHQMQ
/N8/fmKPabZyHsrb+6SO8prTXLQDRisDXlbhXmX1wYNvc6HP0IpsCdy+94jDmLIA85Rm8iL9Zhol
StuepOvRyz4eEkztqPLXMwtj4zzpyNlhlsnzWAWIgSGEN6OxYIEUS2b5Nl6fqbnAPJSXI9NcOjvl
QLQOMYomZly26IskDrQxib581gB6OxSLIOQVKVkU3+wactKD6or7U0hitzXFdITBtkejsIWkakha
5JhQLmbN5ffRa9NlrKuCsnsgR/wc0zSnWc494Vd9VdMaUSSitgYrEI3x6P43TUmAFPM0HcotJqcW
rlT838fWPvMpvf0CzpiwBbGcTR2hWH/eyOMoCdx//6RmfaGwP+fVcWEskKWMFVKRrTdtYZIJl/PX
i9GeOngTwxYEFlqdBMGKLy/Q7YugaYuoSwPpva4b2V1ETo3J0ksFnbN7g/rfiDj7W2Qhu5kw1ttB
3qvwjcIX4ZnwFVU7ks+yWMeodjtsZGwyxTlldkNZJLv+6igSbxhNfLmCZ76uKL9jTrxOqWQSg+vv
Z0Iv5pk4rQwl5rll07GRdPxPLg5K1POVI9uF7StllQgzdYoOK/nw811lEFEzcwpD8E7dWibf+iRU
v9SE3HS4TAb9Vytio0rbflRZCEiFXT8/CDXeXvq/4edc2MvH8juUD1qdvucHG0zXnGL6YHzUTgju
S99KHQaIpu+STEPMgHyhdFUlggAIdkWjlMCN9tghjpwi6/Sg0l4O+2uEcOvPM4e+QgemmL/GYYUW
zrmDLQCU1nn4laEO4XNXVU3a1rbsOIDAD0fD1gQYD057lLgOn5SE4Uz+JG6mpvizDm64Zk0VvTw6
hfvB5OuRfr9/mXvrOqCdcqTOYv6R9e/M+FD9I7k5HJ4J7OO+rbYV56dDLdqFBlmakAbXvcoGh68u
AIeLYkn/iKCXeOUJXfQU6H/C6QLHURt+tUxQKr8+67X+3PXB+J7wIj9ioTPs5UoCIt/jVJXwkAcp
eCMTMpwqcBEjMrFROSvpxZ9kEhePJ1JekMdFPgP+AmxjOaoK0EqCcww3k9xq0P+/UFEd8T656BBJ
VVx/2VQIaeVRH9uSM1/A00ANFJ7gnrddQBrsKUipp8gaPPwPPce/Z3u/tMC8VOktLUCUj1ge6/oU
DIH+7DuYH0FxgZ2q6YoGkwmx+Do//5MCcDQYIUCG9Kom65IjIC6Nm2zFb7/qXVOr1t0V4O4bEky/
kHzmojBaqb1FuQMGheFpZ7ds7ZbM50tzOr0Vqz7PrQuyoyGeu1TQvofWd1UndGuew6jcbP8nAySD
HjoDrAsFxd6tU6Ox3oOCNVseh9cAj8R6zQUXimFBts8p2L+oXdo5A9y9u/Os6biyUHF8P5azzbWY
hgE6dGVBiZhXeDUkaPVeLhQSgVbyM1soXg8yrYATN/NGGw4aV+pxgXCy1QaWcX6hU3jGevFohy3U
P6KfI0Hw1Bq0RTlBjDxS9sDOydfsP9mk6yNhv9lzpNsCrer9y9feeRHgcA35upypfclYky1cpiXm
ubj6l4BV8QCKzjXQltuSYLZE9jRBSFwQ768tXboT+LhWq8CfQKcfz1favZR0gjIKCzfPBuevlagE
Kz/NPhNScLBmls61WMt/ufvjMYeTEiY2nT5R8CbMbmhHa1Yk+M4dC3/+9vKHNBA2hePjMkM3O/AU
E+SldusmxFpIcvocY31scKNy2u+b1R9ugAvRaO6yPJF3rZ8Qd5Hlb47fREAlG/Pn9pgOfzudwRtw
I/wXrYe7vrUraJYSNLHYaBJTXrcIdxgNzvxldky1hJ0WWknCNOUT2cD1CfqfOk2bH/9wJ9sf6vA2
Jc1SSzDnKGzMrc4kxwmMCaQcP3Y6MbWAgbPtrnrmSscuk6tnYiKFZPfDVmQHOcKBHsyqm8f7KQTx
EKpH+4XO5yOhipGhrK4Zk5gZoGwJpksWRbMKemeBNwJb9yulF/v0bjvMINIWGthsIhKXf1dqOAPR
O3XMoEwcXFJClSOIdZKVZ1c4UvWuL6wy150zsY/xbvnk8rMpgSxbrSBg3A9TvgC8FTlktsGDXH4i
SN94mDjF9Uie2JYU4KyV3YpHrFbNWwiD6+I7H85k5T7S14fYE6TF8OQi9dh/uYdfdvueYvmg33qQ
KfqDnE4/oK8qnnW0jn/YuPYNsZAPYNtERPnQmsovm6kHorT9iRbmRd3KCLq5RXcD2OLepAFGrS89
ESHMNvDOWl4yXQKDRVvkEbs+GOsyjvUEwl4dneSxLTZy3wDxgb1dpNGNUr0J6znv6IPuv6lyPP5a
9NUsl5aAhQEs0FtB40k8Mbv5NX3DCfPp1HBA2XqvXWfzScv/sFHD9DiJGEs65TCQgsFh2qELJs9h
J70kjKxtbzKf302aQu8dpKcm+vrGbRoCtKuMVV4IMQKeqvYMGlfdmkGzwy/rJ3M6Fbj5sF0r9taA
RuSh3ou9YeeDLvBdlZcpbKMOU2X10sIt+abWz0u/i8ljWC8faQbErDXYJED2oWApgktWKRV5Yktz
BA5HucqXsEY00k5jwkawqvo885nGYdy0u1sSMPVsMO4SpC5G2wt7l89OgDX3EL0kjw/QAZOcLRE5
DDaXXOe8qbuAr3zMmr3VZiFmnKzewtKJsftF2diW+YPbRIwj7nbTqInt8tJi1RQDMyoygfBMe7C6
/xpC8p0W7So4cedXoBE2QfSgbnrXtdD5SXbOIotQzrBVuDPJnUKFBnOEPdnQAFrDGiy9FioVf1Oy
8nhaPuXHRtvpDRxtjshSyhu1MgTr/LXuQFe6CyuGy455k8RWwiW+U7nogfhc8Cx/WOg/+K3gZXZF
2pbjod6d22ER6ymT/RJmFB70+30fERSdZhwHOOg/EZ8H6AO61LWXDnI+bv8cw2W0M0G2h0Z1OBnF
mvQMRSrG9k1GyO464Av/yxIO9I+pg49Rdyi1b5hUXKSDwVzvVZODfjF3a2Nv4O1CJQ2klo20Vcc3
pGny+lkf8B8gVLHqAl8BI7rn0t1YLat0Am4RsJZ4KCaJbyji3il49gnb/ltzg0oi0XylhREinjne
sXEGskfClOjTEeK02E9SoWcEwu2KI0vN/MBvKycZDRm+I4fZjNzmtyZUp4ldCLudg+oBqqOTxAK7
I4J9yo+w9brPMIeHXCVB16JGbDGZA9qgvyLMoy22GyaPWRpYrmFnCGohvvTEl+1LrgnluCSsYDth
KXRUrFB+Qn8vgEQW8AEYl0LLtxMwAojVAWyoGIFn7ESbD7OQzW1x/RfQDtEFNq7HkMOpNlLITRVw
XX8Qd0nKSnD9BgEkKwlc4IUS3j6wy1bz44GdEYjeBeC2SYcSe0peku1u23ITi01AuQ0rLTD6iUus
78m6FJm9y15fuJAADsVJqMd13q5HjcG2pAekZnoYjnD4+EWx8JAoD9L68HGnCHpG7DseHtCmFixW
PCwUeEcznKXf0WCeLyEjcVW2Dxc82I1384mlGGrXzfHZHmSk2gK0nvLCz98wsnBG4rqwd6VaD1Bk
UoX0eFeSce/a+DwsFMpYTaGx+NfgL8YLiW3briGRjNwDhBbSnxLYpVK4aPTJdLX7g8EuFJ648+sY
kqk5EntO6tSMZPO5a7XBp3rgYxxuGI5UccgjaYxGBBcaF/88is4hluqpE39gpq8N0HfgaV88/jlr
OVCEDOaA5jCdH/oSxkb5m3K0kVAPT/PDeSKQULY5YikW8QEOxumqZ4URwjvQW8tE4FhUG6C42BR6
zgDohMU7inmzT2tTDdp3YixAwIR++NEAObOxfkTjWcN6eEX5MQFHhTFMKdiCChKkZ72HtlCFPSK6
sVNkwmuYcmSLj9UyyYOQvQ78w2Bp9cnK5Yjsjw5edFejwnT6f3AV+41cDbx+XyeeANXbo2PEJ+FT
bOqk1TZbEqM5hdxHUDkOJmJC6x9TLO/HhQdRJ9/tNet64mqox7aRKRKd5SGzLByHbBwVkc2RymWa
f0JkT8xLFub9Vf93Tnf783mz9CVq6wPKnEQxjFN77QSP05/ZQb6EDgcGWmzNeZAgkw8wHGOAzDHr
a5MEy9zSVo607/zhe7B01DB3KmTaYpVHXn7JToh1QQauUdzf2kGcqoSsEXzzg2FcNba36Vt2/Xna
+97UDPcNFGogOeCWcEdK89Oqm7DRrIsZENw4cZGUnKBsNbNQyxTSLGeJhCa7h19CfdDh1fNc63YG
kCOVIZ7LQL62KIui6M1oTCmXJjlGzfeORgUhG4w3BvObU4FkFmStLi5Xg3JPlvaQESOXEJumQhCS
Ck/uH3kXETJ1KobyB/0F3RHfzF7Bxdo6ttDgb1rEH+uM9DMxBy6ygqfCBdrvBuRtTr+6fZ8YG8AV
a55NLmeZkwh0Ve/xC8Ix0CjHXR0kaWCiao2IEsfNBzj7gpO1GJfRPqPJcNCf1plevXJH5ioYxwJM
Iq2pqnhy4hlkJKcwnT/4e6VPx2/hJ7/o9EvO5wKF0YDOwJykomh3ErYa8SLZgg/TnuYuS7g1KsVc
vZ8Sz1zo6leRlOKPs4flAwLrTEBE/aM7oR/iZmC6KQ/fw0cIMrNZ0Bsh/sxkargQw5tPa7+yGsRQ
/BmrHjZ/yMZoqRJfJRzR6YIgsBdNvjK1c8INni/niGfhM1h2agG3QsBARM4R2X/k4LqS1yjWmAsv
0j2yXNlRL+ewMMC54+Tyqx+4dSbHFqSTbxsQajE71uBARBNIfl5iYJid8hUZnojGBfOw+ky8EWLX
S2YAzTPRX3lzwlE2ZS/ThXp4BmCVKy3ACY4pedLw87UljsNDrFg+WzylEI62EWu+Xpq9i5f2yR93
b97eDKprvRsbqEGMt3V8ScOBtN5UQo2mWCd3rLsEKO580uPC3s8q/FOolGFXH6Wikwk88hm/SjdS
agA6t46dIGyW6CMaPHO+Fws/Zh6kaqVUJaS43X18gAbFVDcYhZgWMrpMhfK/QD4K6zkI+YBZLkqo
nawKJDlR/ZrDt6TFrZClupU4f6BTF+vLvjmV+oO8ER5Z9qDqdGADawttWvS9PPve2w4xkE+VHnDs
4KLR04upJABrf2WpDbidzD35eC62JP/iQ/J09iM+H9SAEsDR3cI71xwMDdqaOACrHp6xtsCTQ5ST
RawAg9W9WwjsNmb2Yarx9ebkKHX8RvFEvrVYy5SK/KpF5KFPiDa2GgZO+8X7r6YdawmauuNL50GL
UD5ldk2naNqhQEe8C1KuG4gnF0mTffgx+7Tgg4VEf967OOzaWksM+8kUGG96B3sdphZBKk5sRdG7
PIxWPbLLP+YN8XVHcNxHqdpD8QqQQhj0EHn5gI/xGljSuA24Y7w4Ei7jYLy+7p3wdLWsPmcbbc0g
hYI4sPLSIOm4/8MkxFK53FNpDgoIHWpY4aQUZV7juBFP86PwbD/vIp0SlTbwa52owWJA9vbA6HIw
StwHPa883Ycbi7f5xHGh/2hd0ZHZ5jh84UqXPOgyohIDttA3//JSGakNBMcu5cpZM5mjoE4qTMOt
rEbYxNqAa9Q74cZw6Mxc1nyHgvoHfYoB869bXrRgLDyS8k4s7pGDLWyxCXPjtBmUrZzzBISRRDrq
JQb2BQnPEYe4b6OWApv91mxtUhNjbTAujvIwdul8nIe5GePaycU2SsaJepGlheHba4iX2QZn8qVV
IxReO1LWLZerTCldu10aePPljfK0UcEfSQaZLn7gtxmPmImX+qx1Av4VuOj5s05ytEZroxs3CiNH
KrenlbTaIP9Xwk+DZpmqWoIGqVj1ANBLwk7EtZarfUMaMykv8f0SrpWoV8Jae0sroXu+IJH4V4sx
g3wXisQELXwAiWvUFyzoq7ByZOp3HHOu4DcvonV7+Y9hV/tmlEJI+VpxFIYk1fUOSyorwGUimpBB
nEZ7gv1fb4inzO1g+t+tVG3Qv1d7rRnRsJx394Qdd2ABQIi6Mc3QMjjpIlWL5LNwJ5BVrLNtmqzB
1Avzvn8VWgSieXa12IsrvmECIUeH+uC9/aJZnRpIHgMgfkRvqEv67piO0Vzskfls8OEiV/biqf76
X3YPkWv/FgwcB8GLjzRcn7MINzumIJA1nC+Kg5nHj3/LfYmBxGPBCgYHys9FA8SDDVOV6UjITR65
DIWIpYFJnbJsCowS4j5EsnnTL+tvuvGswE8yzXtMLarvbKfdurfbKtQh0nuKzvFkm1xL2MqirZQ1
/c5GY4E1d4LWl73nc1eYid8Qigwq1MKV8UM7Cy8eZVHEe+PQ38XMTy25EKhfKDxduwLIVgQZ//ky
73Vj4QY+y82Qsf0IDsXeuEK9mSOIRk41gneOTI1iGpZjtlo+CMAFL6772bUUNiXSwH0EbM1oBLke
Lufes6O7ZtM1OUriU0BFdGzpOOPqXA762rTlmPniw49yFeFNn/U17hKLMroA/zWhjWMFu+7HtZzW
BPHuq6VwJzHs2aG0lss6kQhfUg6Xn2TYFN+ZVL5kNwFhXb7m12s9gBYgoytuwQjCJyrEQKg7sgiv
06/VKWgpb/WDTfIs10iQfo55sryyIgNx5bLJ8bdprv+a4T7UrsB8P6waTSs7cp7FIs+uLuS9IBUT
WE8rJtiWGNEKz43B+cvxXwG0/ewc8v8bvz0sr3ClY/O4ICtOrR5ePg0bZvq4WAoZ0/Ptc844fMRW
PedQn3FveSmKCY4FDz+O3NMyTSBpzkcFIGpglNcbl2HJVbbzGM3gDwCYHeT4HXoBt7F69+f4bscv
+2jh9NRIeSiX0k+d3uleg+q2J2rBEnpITNdxMjLO77JKuxDyBtXDmgST14leimhbl+KiEo1hkhdT
YLFS16t1OceEcnQRLYpZCDGSGKG6asO6hKHeU+RwTHhg1M8qge7jq+Nz8GcuLh4TT2KdysEbry3l
/jkaSV7MW7pgp5iP87I1z8FyPAn80x9CgtuNimk5sOJOul3V7j1puWPpGwZ0vDCoFlhskOxkwhsI
APPKMxmzRFcC6VixAQYZ9c7WO6ZyzYP9PK0taCftKzEXqXZY+KYM34vFjSSW7GuBJVORJ82iUuoQ
Bx3xPNDdC/La5OhlcA2RnZZokXt2YXoI3UfXuZ95U1U8pcEiIHaPR7CDb7aSqspXwO9z3sAah6kP
RBlKJIvZE5sAWtwcEt+Adt1FoKpbl+6DL39YLCnSOP1TKUurRXaZqmmSQ7coT58ZbP6Gv0vxrmLG
EjHeDKv4IJL0q7aFjxtnORHCpPkRctxx38Uu7Q+IJScw1FnKVDFAo3yK8n5YK8s5bYym7FmAYJ15
sdEMdNfSDHV+omt8uqIyktN1qb67t5uglJp/duTG1Z30hcvn+zke32G9hnh4fqUj17fiP+IuWfuS
C9vYrFU+kIcDGETRao0KcdclT+HpL0+Tti4zsBGJ2dQSQIwfm2aNvsFGxLSIVtBx34MEybELWqrY
7F5OC4uCwS7EPaDQDe2Vwi+zY40tyriarh5xGJlqAgSijnNs8PF71T15cR+BN76Ig/CjeU7S6gsn
eOso7A2bskWVXt62aHvJuSXPzsXBhNM6ec4hRIIiP9Wp0iYt5OFAp/GQ0h/KzqAhvFvyWmQZDX5b
5TEGsIO+hpAzZFXcIqgaabNQal9LIDcr1KQ1DYCkU/HfYY8weYatUU32n/UUyXEz04Z6hoR5xsCr
SIqvV/9gQYlJ7eKmQKBzoWvn/vPEf1UodqJFshFYD7wDPA6juL4hu4RwpeBehMaAdE7VcE9aZXwT
A28R56KuHGNL50KWkRcTEDIB2aUwsyz4D4jiTjx02BX7xjbjrxyFTAo7JLxVD98VTW7bwn/GVK95
meTJXQ900Ub2EPGuiyQ5QBZH+TlyBXeMrBb+Q0KO2ZdSf7wrLSDfjTXKyA5TcpTceF6rFqpkDny9
EyLH/kRKje0cByXLP+bRuLvvejOzTUEW952oBEN9lW0jPgaza8YS9RrbdzERxiPC3KA8HbN3tyPD
7DaW7NLnk1WtN/g/IerTXhNeoxZ00VZYsSpxltG6sjvgpAagtXNWzMhoL8S22VjoCx1EVuZlW+qJ
7ViwuhjQusiwkkM25vk3xWJuSjzLVSNyXHs35bm4ol3UfuE05qY3dqZub7RFB0BPZSEelONAElj1
/ssSmhHenOWhiPYreaJbCNCZGav/UdQEqUNwaYMvgZbVkSgpExxRb0gs2ZV+GSRYVY68O8skZFcx
xhCXL+fsmQgFAW/PtHQwJGR+ROZz9jy8M3lzSwpVIhyI/fqNQE264FGc40Td/PBuZ2TQYZNFwrpf
xu0xSbBRcTPq4bvPZhKASlV4m5T53b0V9h40ERUuNYcwCmBBOkYtk9r9SdQjTMM5j7M13XIaBSNV
KdqhvoWfYjbSOtuhrl1mYXDKlMxnZVDDzRbUrIysOyEj4Y+Z92Tv2lCpIyxTV1UJL5AZjpYykV4B
ShmU9QZkDsXoEvx5DTFHn7Ru+MniireomTbEnGyw3nKrBQTO2obttIVJqgrTK5Fd4nf7B3L73Y/e
cRX+PCbbnAuKgeOxoPea6ukmOpzL/PFsBB+tMxmNqzbZlrvokrLBJiLcsujosV4UF8Cb/LG/TkUp
Zgunk+UaM/IcHPLRtV9a+7AGD/AGOucpQWSLIZSow9D/b2Uv8GKa4xdW4Ab8aj4pdNRp52C0BoOo
epiv5/eFYVUEef0PCPCnLt5ZNNca7a9hMa9YWLAmaBj9dekULwkiKMUur2vvyaYgUgx8WdQ7RpPp
ZraynlosvggTIqabblUTijZlVtZwAsyED/JfMCjuG5mZ8WbedrMabMawhdnljOWAzFZG7HPiLUjA
jCKoQFONf5JUFY6QV9PreHPA/qN+O+9qMpFrqwZ+g0RJ+ttk2vkA/TzF2Lt3OX1E/GqQp19Ntg5e
qE1wKtyr7bOcbtdm08TA1Z2GVUOSUjKLGepjspI+ox25bJtZ/gmg44rlYu3wZvIiWU0vwDtOm9BK
+H7IJXTPEvV25yEPCcZD9FdN1PguMUNYXaN7ADCeuh4Taiat8wX/6aZVgEq/TK1l9x8V8+gjAQnW
Gq/Dsqqcj3eJVvDUZ1naT/3Nk3vUbk436RC8clUb6bhTTiLaRQyxWIcX2kYOZENwkqpHI5R5Xw3c
REQAPF81pG854X9s7Zjj8fyg3wv4/fW6b7fth8AB0U8ibTGL+rGqhdAAd71zLBuDN/CY5ob3wt8F
xZixGXvkH2j6oyv5Sr2yapVkJeI2XsCmY62IEbiEWw3CfIN6FS0J8KadWICxxgmnHUHbAnoTFgw7
KyDTKgnaMdvnhxPAceweFFBA9C+kNBYBdhgJQthcVJMla8Kc0PqoKP5s65EAd2JypjUr3M1M7DE7
qO9jFjeYr5JE4X9Pnm0UWPnczfE9avPTzbghYiApBn4S8rfJ0L2c9qV+wdu29qv5TDeMPdF1WSiT
VpbEHQ4zqlwh/gGbF6rKy57D1Ai/25aOB9o4wzcOdW2AcgFsJb7nGvTUpol74+CH4Y2oEEPjh+Yu
+Obs7MvxTnkVqHV6z1hrCUVzxwpALtNGcedrPm80x2nVTlWpk6WStjyhFj2fpY1/5s6nhD4KV5Lc
udE5wWTOygKT+i8Nwxohib1bgzIrnd1499tJJeOvbNXMPjTwkkG2x8gGv2Cc1Ayn6xbuWpZ6P+5g
mBu9ipuQs1i80WPjkGShOheUdG8L3X9JIvbBpHmdPNiRSNtyq+zVT3vFT3AmVR9pD0xb6rjMxRDF
JWjpXaJUcd88Rfl2v150F3Si6w2iijGpuTBuksj7gP7zdb6xA05N1Y1Uzz3qAQ1g2CrtCibSDi0Q
NU7+OKAEraa6KH1HggEGp9EWLZuoB2ZyoUb2Qn1eVZTvEDlvQYHwpmhgLJMyygglnQx9V9k5Ar+c
kbW9NlgHRGOHfaFNYqEVx54sLMucSRXpXZsTf9gxIJNtS8IsanCo13QJRz+DFtRF3kfuE8drf1Jc
SVfluGGfiyUxLLOl3PLAgqOhBlQA+Vsn3IM9rAed2PA2I8CJ89Wwg4GBZK0ITp31e15yPjWklzHS
3iARpCJBW4fa8by/eongNeUlmztIcQxuR5uJRs57ed5DicdlMnpcciljOONPeR11XexK3m51cYoE
nwfjO22UznmU9gf8QIySx2JNioTFtBlQprhwKUzSk7vXoBc+3g8WAdkveCQZa8HEOKSvyBNxYxFR
VP3MRP7agA/E2GuCictEiGmTojHU3EmezpmxYYe0YhnWst57Fkqbf0G69euNXILJYzyn8K2NuvO7
WBtZH/oVlNa9sTHK/qsban/aXlPV8I5//1p74yXKrROqHKdtWvXzJeRaZXhgBLGWPrxM+gsyyixa
P+G67w//ZmUoKwFPOTGxT/a1Mzq+rKap28PzqvgTmmcfdOMLbcObWQU28y+Xa7171N/ANLS/RU/v
HI7AkR8nBjs03F8L8AceLjnWQS8eeRSBy1K+BE/WT8D8Vt1w2250ikvCSnyTicLu3eAw9ScYZ6gF
rX//r2RDQvM2GPWGmE8W/lrVL7+uga/uMRf4pF5+xzqwZKBbUZ1gjZmIYBvbklcEjQVoGPOFZLe8
7dMn0HhF4Fq7AfO3r15faf+Z6VkwVJ8AtvxYTTUi7J+h4/5EUzAu7NhpSG821nEQqfsGacKjH8zu
znAMgJZwkQ2zsMnYeIUCVBOPyaJGxZyTWrBU4yuGPNrVRhQepMNmNtv2aZTGtQgMqOMFYXo5/zrP
rIBhZkb7OLSz777OruSVMbGTCjRwumWpcAGcegyQyradbHY5VPJXk7lu0Tf5HpgiY1BnvYcv1GcW
XexwEnMgGT0ik1R9mSARfjcLJAZCQSwOXqABWitRfP7hkRQnucRPuIIORsjKQD/DfDwv+Wd8Xupv
yAxPQGsYqjXlftwSy9fZvRGWSoPRO3hQNIbZReKhrbifBd24I7ckQGwgzC0VGt4dRogblNWjwVX6
ACS0D9RXXSzqrl1o3m42h38G2/LEvZHn/YliAZFsmGDnP8hZlN/Cd2P91+TNnd8zcCbR0FafDzvx
gDZdtQUpePNHxgJfoM5Hzvzf6RVn6r2QDJlsypbSPHOJJaU6rj4jGbiTZI7SIRpkjiaK6+2aBPtf
UIZWY8kHF4x0dF/bb/WB/JRDtBDrxmiE3tjeVW/uezidnQZwJwDUg5j4XSuBNnR5aFlihwnyIDyy
6kzs5Pj+f9a8Im7XzhphVV2FRwiR9zyv7ej9w79FtZjPHCwPZTN5CMrnh4nw7Vn0iuBXSyDCyxoR
aUo5oyvqfs5oxbybAKETH6ebXyal9nd96pdznbherD4vc6XOa1EEW07U9JJ+VIYqnhlxcugHKydS
ltJvm/0Qv3lHQTwF4XqthZrqQSZJetQyJYOwVYOSh3562NNgX71I8z8l+pZNcHaVftmrmjLcZ28S
dhpkYJc7/+n3rFxevkJ+bYqtILq8mutt22V+2QUgJDRMigeIcB2849S2+89DRnM0qhWy/AeqzRIr
JrIK1Frqj1uEjSui8TQDquLz/liVOhXZa8l2jZa4OBpIKP20aDWiajnTT82B9nS+tx4kGljXaWX4
V50MB2BAOfVIRNKFjlGoF8BvATDM28yRaod7A7pewsyaGbojKp5szzq3rBQulsEXnYUyi9j8hs9C
9R0GfPyxXD1GFVsSGsz0aA+80GrCfYvO+vfosVNZtGp7UBtLCtGzXM5p2ye1o8qfhhLYRDLoSt7D
lorFrp5dVCXDAleOTVBR/lWvVHiYsoO4ThO2DnIVq/YTAggDq8HUBIEIbCHSUgPeh39X2r156foW
G7UPJBoxJJ+QCC5MnYskh8SuVmIR9lOJyxGwNk2RyIC3+doR+FDuP+BbmBfajTexuey8mnOvQ8st
BbNMCbpj+NyKsR0iuq3XWlLqqovsYTBRaS14Ae83sA/5ZNX/z86bPXJ5BldDI/dK4hz9Vjvlckji
pOhmWYE124fFaU0ZXWL3CcxDRlED7Qxg1wYrsJbZiHV2PhlLGtS793z9gw4pnMZMEAwmtHGcHJoo
0BRRPtiWPyMtufXsQz7yyPYe0MShumdagmTUSVfc2ydI22qsd7Jqjj/U7jvDK0fOC+umjTdox6xQ
mn57gT8hVP9IvWusPqmGLW5IGlhPN2CiPALV58m6U46IV8qakdbM8T1HMFNYw/PkBaAXU7NZUIia
1g3mPZOCcM0hrZwTX5Xz2Zv62SKr4SjKTDPZhE/g1TW0FGa8AoV60eoGDpGcMRwy7ymAzEQSviI7
cELmQkA5VLQm1keEQCAzGPUD8R/JVqeDmpYNeRQOnBPrqNTMyMFOZivP6g0v/4X0Ag6PLagQqyxx
XSgiDJp/ZZ5nnfRrAw8d5zQOmm/J1LsftXsRAUi4GaGIapKF9Vu77S3+rEwbYZ3DLqIaj+EQv1Za
H/goKv+dzAgwZdtOukx9TmXjIZcEj0xz7mTlbnLqHNjuWnrLt/H4k3r16SD93sfJ89wCpqGLnWh5
ZLgeITGbYtarPMsvyndCaJ3uSifE6vupHJj+nxs9SbMpy2+EdFmNXcftGH8BUVZaJmi2QSbHJ05b
lSRt30gzgzY+kJrNeIHixXmmZJdBkCcbv+6DlUHOYQ9Brct+lH7u4vLu1Go8VH+VBowfrm9cAQKu
hUW2sX194GoNTzfhIWqEyH5oyG8whCaT8unhQJKvvG1c4rMIVsD1wA922UcCOfC5Gcx1JN480WDs
Kso/B8ji6m83KmLcMAoO9U1I5i5QAr3jl9A03PutUEOWMewK7yus6xdcK080qmmAysNXs5foCVFe
lhk4NDiWC7W/CjGvvXvDJCjQRaBH/yULahw9uZmu81pmLGLVfewlROrmSsapb7II14MDov80N4D8
aW4knm6m1Qa8pVoGCWCvJ263xMKAxNf1tJk9wz9i9AEZc4ZEHxFZkA6OhNKQQwTcvlDk4+EyR91P
WvEwwU6EToYPKmuEi2l/eXCSWbmfcrUpxxBDFjhk4T7Ib6ZMAhiIFkfZgHVCd2dfsQh8EPHnkYE4
h8spbrGEGxAeevjlHt1E1O8qTcLijJdQQH9Lml1lNkJhvA+A+7Y2Stbl6unEqgLk8RSRJkcoemVg
at+CRZNiscapNghMozVgcMvXXPthpZQ9wRjdytRcaRSK1vho4ugkZGD4mUXmMDITq/hYM+H5sbZJ
GIgbB47XpCR2glSChcdyq2DYDZXdc5l9mWFIDt6kBM9RLDq+M+P/t2TAYm4UmJY4GQnnLO/TQVck
QPiA26ElKlAoJl29EIMgWmFVe0VGZLJsOa/rRRBHZ9pjU6rlPpb7AILDbuVDcGLPPyLU9Ms3BJHm
9lhaz5zKf51HGOiTeAZLTofRNS8VDoSd4Y+Wc+qeuVvPyxdddNKqw0bzzoDeS5Mi5WNerA7VosP/
UCp5OX1F77Bz+z4YHkr6kIFJCS+ZSThjp/j8l1c28S5QNUVCCNqYp8/aGb2Fq+92rxcgI45nySh+
iJRydVuhH4TKGhjtcjrSpXX+vEG/sMBhh35ZRh77FtwPgnPb5n3UX/5atSx3MXYlYeYx/3St9BMR
Ipg03BXfc5y+0UwKnJUkfQdTycquOMfFkWUwmldBLUWdao9BQ8ay4TMVIN/LHPo8TXE1wsQvdGgN
uD+3M0QgjPBNpNnVL1miapEBBpHBlC/sycbuYi6keQWSQxbtXuSOlb/gAO/+Lk7czaUjz4Ofyy0G
0jAVg2HnBha87Xwx04COUAAq3/HTmGdH9n+QNrZW1PGklv1r8lYHiAUEr/xFfGtGLYuz2fPIrbQ3
VXi8m07txd1IeyYMZ2VFLtIoVUh0uaEIGyrxY2whHk7vB+t0958I44U+ioyIhGEPPQ4cByE6Iz91
QNyF4EWdOTDBkb8WDqotieamf0swt08fQOXxezuuWaLY/99b1XAZ2a29MxsvrLwjQ6Ax4PkDNJXg
nH8Y51J2gh+BoMp6135qAZGggqFePRhyqAPivJhv1Zb86UNlX+M+274UXQG7wGfUp2o+LOIT++Tt
u0p9pJUSSZJw8/wDzeb/OIJs7N278WquklnilBUnSLsfv9xGaZNwU21xyX0ZvRoqqf9Fzj1rZcBh
TET4NHUJCJZs/yIgZgyyORHc1J+GlJVs1hoMJJfzwVrONbNIPAjgbjGuhBklUyUQVDdqKWrCA9oO
IjgypXykqJk02+N1fUCQME/i510XPxuuOrFi0jPqc3BbP2Li8w+GYDRXF5Uq/bJcGbvN2Varhov7
zr+dLvPp+DvUi8pvL0u8FdhvczZQZ6/Dpa2lEO79fqYoyhH+rIz1NgLDdyWiALBu60GPCVJi6ga1
0HdMhxnEHlsWJAYZTzq+/aOnzzH7mPHDnCPSz9JIVVqBIUBOc2zMhTKv797+cwqBbGp8IIe5CzMc
Bqy95rPCrEqeRbOeX3Jul4MIXLFP14DCxQ+47kZZHd4aoiZzWj4eCd/WwF0TLp5Iz2QVXLUuXo5j
DLTj8AwLlOIb/unGDalF3rVWlNs6qITYWdV07Xh7lC0Y8qiLP8+7+2g7AvizCOkAttV2MQrlMvrz
ogmCyH7i46+RjIqE5NlRZxIUwm16RRjzGfYWRISjnBMiDftwl6S54cS44AHnNZUHsvs5p1ZWRj1/
8knDg5l2fixTBY1PFk9NwcC1TqbXbxxXCZSV/bnQEspMQxor5ycn46W5viisjfWqnibX8C9z9ULF
qJtYxT/lX19v+oi00GuI1EIssVAuZGCajcydWA8fTI7BSMaIjU7Q3CZLU+SRDVWYLf4oerXpG86b
uBXk1usamc4QolwxPFADJCD3hCy+GvWRj+hTnyVAsXb163FirEPa7T+J7eLzt5RB48+x9mJyeGBq
ngMPR1Tq4X124zcOraLpZEeRM2HnOXbdZQZa2nF7iEXLgxSQvnvczAt14PjeZy00vqwR/TVCPlcl
oWVpNA1yNeglcgvt3mwsmTwvbNxaxcTxmEeWnBkmJG6leHqdcDkkwrC3pxgYi14f3elz3XfK2kYb
FHK46gI+tX6kUtIgIQ5jxe+IZw4CCiFdSMReXhWM9an7JxcQKTeCdNUzWp/ybzpscAPH76N4nVhU
Ez1iPQJxnYKogbmZFKV6Fa/8/JfCASz2zOjE4HwSCZlAu7Djmr+0NlRdUSRyeK8N40Ij/PFxLQlG
cuxwb5XsBd8I81L+JaZ1AZvYqphYkhZSdRCJyrDRVshW3jrHKb56rs1NBwC1AgqsrjEsMMnAArjN
ak7b1j77u2KvAJgdfrDhKKoFI75ZjHjOyHgVgTd0PoYD+OUlKuNjU64feX5EIwa3hbFH7JgzNQON
lm1L+9ePjQETS3vL5/y70gmyweiIgybPYocyPBbx9SwXD9rgVFqnV/REkw8L3bfShIgURXUm+SCa
lBOtBF7m9Es51VNkVH4R3dX/waUTszcslj23mi4g7VB0jR5kdNbBwmbIA2AIh6BOkaKzIQ/SEGUC
LaAIMyMEzd30zthGe6wKY6glHEaPWJG55gpsBdNT+4XOCoBuwxAj3J6CIFCwOft9i7KX5AZU0tpt
RP+4/wFMxvWekujd+HPmezaVKHpcXZlkeHBkQEYoCTEtTLqoe46f6KzPiTQlAUcJbzKNt4fEQHa5
m4c38dYD31dPX15g27cO1Iz2KjhAhe3hmMddb1yVtSvInrCbYFdO2/tSnwjhiqz7ufqz+kCOLxmU
QDFEzuTRqKRgDk8TQAl+xYDmkHrsKbxcT6yVGdz82R5MTrHiVDmEBUr/mGJ1kwX/U2UEzrzj903t
deSkxybKNrEIIIis1No6swSMYUJkMA52N8tpI/gXdIDFmWbHJusMh/EaMmi3CfktxXnVZ67vF9A8
Jv0K7C84WDciOG5W/ghZ5fJvE6FL7O289GoR6kiXV0PS+vM5cTcHA/nfeVr31DhdplsEaz75vnWu
suP2xJyRIQrd4rhG/1jQ5U6sgFKJytQAvldinAa8+D+oxF+IILWp17JUmemrE66W9e6WZQk9qDht
oCQfcgNX8sxiag04ivPNNRgYVJDOuH3RQ95rLTBCC30lirfWbTwiU6uz0nP7JUv35FzLygfaIUKW
c0JxQ2tqV/vVBwRioQP7RIiEek1D/7CYMavIe2tKClKU1UZwn3B8h+YW5i2c1AZQAkQKWSPKwHXD
SItexjQNX69Pm93B772YLr2puwwv3qRj+JtoUB0CjK6MJdT1cYjf0EAnWNmQpGcsvO9wZR136U7d
hRD5cwaWz93NDm2+slSmutiylPutaa9b2ZAfFH7VKMLwXwrLhTY0AuYTsGOgrBFYMn2O25xlBw2u
HmHm6fu4mWrGp7QCvZoDGBjGiO0nPoA2meZUgSeAhQH9BMuxCC8O9/7nYLoF6239mP0Tvz5KU1lh
55doVV29XP/vbB5+2JrNWeGKItwQa2e709381Fd4GusLMd83EWlQGbFn8mMdtrKdVLZwpgzfgq98
wvthgk1kzDWZqkcWo5vNWz1NUZXhTqxriT4xaoIJ8hXUpjy75bAUDhQppoz0Ui9p9rdKrKubhQgK
96TP3+l3ey8IzpZXCj3PGkmEZZ2++bdVFaEkTQNvJxX5gFA7sgN4VN/qo13xhbiE9FnOD/ci8xvE
jJb0Ffda0UGsJMpLcAQd4POzRVcO6Dzk+/LqIm/g3KciaoVoKQzNbWqAFm4BdGVt0fZ2f4sgjTya
7ehd2ZoFpcqGabCq7v3N8MrIauAEYOM5p3hYTipi2GqrL55frdfBlv1qAyqhSTn9TeZN4pPY4DNT
FcINYdBeweTOGOTM5xGjlooeSDggP+FmA0h7awYxzz0GZwPPzoWkTwAx61s+Wc+yuUkEabU5qPf2
V4m6nGwVGyS7K3m3R7iC9hUKQNhzdTLsrsk4AShepqAyCBDW9JURPX8CdFHSydG3nUqqziEpSkvC
XxXY+D2xF4xaXDOanEn6KJcqgmWtSPJ9wpygMGR7o5cGkOrMHBIRhoS70lvAwEI4NLNwpbQcyCJb
ZHG3nC4N/g2MCBu8SUiE1bhGq72YBW7Uz3GT2nubNzJHcxhsEOKYvYqzdOBZZIlR1M2V3D2en0h+
Ps1a1ahc5QLx1QjA+YhOXcjVCptEVMFyi5lWMI2VbiO+AJSTEk/80yDK43v2EtdualLdU2l1Aq15
CL26WeM2G9d6KgPbooaET/V7UeJpyXQPw2JJZp4E9oWJ1kNmuOagbI6d4zpE9Hp66hLQAndmaoEi
ADiPlEpI5L2FGBVK6PanwGvH8Ko7to34s7GRDJp1KCND9V9xscZD2UHH48uDxnJIHtLTu6mCTOEJ
ojEoK9yrTJVrczlaz/wUf3N7jfUQo0kB34QJfm2hc4Yao3Sxh4h/DJde4U5y5dT7Re5X7QXUKNLu
Z2UVUAV92HaxyO8zxGJYppqJKRVZMdiCwcC823EhVemwoNMTddsHbxn84nHAWF/s5Rpe2Y9CC9Vq
9l7YGzuLfPwmFhqhxiv1msDdnpqHybmVgV8v5f1WoOisJhOof98UflkiPYp4lo4Jnrh+lEN/NVOU
UrNrDSLjeFEkblA3NziANKQl1m6HURWEunZCUkeFcHhQAzuKfwXIxSlb9bRIvy7PM4QF1DTe6htc
T2pst1xhgDnL1rHt+d0DOKkhsGrnp1BZnw/19ILwsR06JmBwL3x1+p4pxONhSexLMJj8XExinAtC
sJ74QBZ0VyAd1o3rxPTw4kNvQPpuCRVe8R5U7PsVyF/1AxxvB5vF6gFEdn5ewSNasNYrd9+XHsxW
JRTMlA5U9E6k4H8PsJ/6V6dE2PN2rFr3HK4cAhTVEdo254Fixj74Mb/MNCBjOm2xoNK1u2jgiixo
dKdzW8CycuFnqX2YDz0W10HohQk4095L5OM4Ny35LksyD8XG98yGuiHkiK4Z+A7/AzpHjTH5cKYA
PFJfGBAnRgClym5MnRY+jcVZ5V/TZhzm3WgZNk4zbr0DaehJruhvBqFN4RW7R98pXkDv+hRPkQSz
hpwdX+soY12KpNiXQqYm+83c9VoHXNWv4hAumPH99B+7oSPlEoQWF80yO7pr5o4K1C2JH7SnKqGl
Hd6YfOmvAWx0/hJ2Psc3tB0HXUaGvsl3IN4yqOk5rAoqywBCdUZ6a4Jfs7HD75TjnWAz38/zcrxx
LKsrbSAkI8ZZ75rzzNSvwAyeis0+c6JRS+yTO+yawYehrIy2KFqM3lVKVkXRekL95kN3mjGK7faI
Lg3xOHFJsYl2vsYLtPFbEB6JrCkV9nTxo9mCSrp2ymeaSwEuK/Jr9h9x8Xqi7tOUjzu1meyfU4qs
2DlEsELg4axWEEHHjr76r9ulCFx7bbMHZsjyv1ADnSBWWrW0/9rDFc7qyqe82hDjujuj1bGtVfl7
7qMtZG1V7faa0/lqRdnASvk5SUYUNiV2yHHtmUr2KoyJDTUQ0655Pes0K8kadBoHp5dQr3jp2F7N
iR95VMuhRBj5nN3U7zhm/gxYrXhbFHDF/+1JRK8cDJqwNhcAKrp9Bpx6VSpF4GkVqLkQLLy3swg+
8Nc4YIxlqcdhwetNZDr3icAWcypw2EBUwbmCqox1i/dKo6QWTt0Ve3VR+A1eapBUks08+66vW0Nh
/NUh4virXz+RrYVzxOkqTe7I33W1WKnfl7mC3kRbHn0OzElWSX7ByMC3tjmjRqCQYU3GMzAeoiBk
tgks3EzG2KOUjAouve3N0meSYwz4f0wjP6dKRTuxbdk670/jb1UNLADOqCeOH7A0eWWKCYtOyBMq
YV/nyAiW2MvpDfSrnta4kc+0e06Fwbwi0am+//GdjwLrSmAvEq9HvbN404qb4XDoWGRqO/NLn8j8
dJL7tUGER0PAeF04OPhjHcgfbOjl4Fa17MYT0TvSzmLbLnt67bYMMNcikqtZLOgB+wKtGF2KjvT9
4p9FFVQaFeaZBFuJEdjtbYHLGFYTP7apSms+s0FW+xG7ZMbfrhX4Z985r3E70sY0SWw6C2CJoNOV
L2X7jfeeVeStO1jsKFbqBJE+oMWBtgoPaf+wDXW1ysTDFQ86DhKDf2M4A/uJ0AqpNMKD6jNNLr79
/3E6/ITjafBoNePfoQXzu2Kt2tCmw83IfD4WRxWh6G+ibIDmQ4ac5/MnSDHhVUKRt44At5Y3gcui
I0yD7Je41UIFLxArfWjc9vH4T2yobFyJXPP4uL2dBMMPdcxXzf7NG34vMmr9dKoxB+1xfEkaHAKe
QMFSfmvg2MaeI/tDgPCwWTcXuE9hIo1EIhfQFMr0bovqe+4JXQD5/7QvhVgAajYspslKZ3/QsJGd
wFYaF9uwIBqGYSCSrz4XafgLDl5fiUvMYjy+NVlpekTOdgDcsFgDkQjmCokk9YecVeDy2dWpADW+
f2EVvvQkebFC3DOkYb8R8Yn0DCg8RqJS3YKZMGQngVLcexsKOQQBtiIDwX4vEbYhwPp/OXkdmN8r
wdG7eQDaIxXohDquRlh9Akdwk5ucLEk6QqM2v99bqcFtfs4k5yeTrvZUf6aJQsMh1TNG7IaeFLkS
tJ6E64vpviqwgmZhYVSfUP2+CatGkLn2hYR3pHtXjB8zd8W29PM5tH2vysN0kDr1fevzWOgoZ6eW
le4yrD+BnIo/F6j6gRary9Ie0FV2gyw23cIOkKtEh98nhW9e6lkb/QZdihFvtc6ZxGxcYmtK+zC8
MK2sXhX6sjGLx9MghpyawYYeukaz3rsn2kHiWHY+g3ABEDvuVBxVbgUFGP8g9lfXI6PNipndijba
XJRK9LtPKlMlKa0HQ+yvH1KKwatIe6LEX/NU4xei1qIHoA/RJOJwzBrHRwecMxiX01yQXFuyHLWH
NgD+RTCg0pXFuJWuBtX2FraGMoCoqTbv87x9Vp69hVLi6hHqzzRH0S463khxMP75U6syn9203ji5
q+MSjAusuhc89gVV8yhvs1veLm1vOouTtPAlwSuBeEDw7xI9tZkY9Irw/fX7rNkYfcMi+Q21Cgxn
d+0Kx2LqimY25Of1BoSNERqFP/M+7hXC/Cd8oxQiDv2DyFyKQuluqgsHn65urO+/6fh2NuBNfpZz
JnTgKhvrzBb3ja2l9WYhnp8gTWVr8E7owaznGx0Wu+fNpd9Fen88ZEoMdddf62dGlnz4svNCv99a
SIvji9RK3wT7N7GvpYf4qu+VYJN7UDaxcvHhkvGj5Xt4XQ5X/Q4WKaU/ziQEySnwxF4Sp7qYP/kl
xQHLKPT9nRAbnI1duSj9aYUvD4UOIoq+wci3MqA2Oz2qaBISRDV7bxFp9VJjaxDkMLQZG7ucL+we
8O8NlKfMDNuH9cSmLk0aEXpiefMPuyNfRTz8U9ywoLvpaT4H3xNAOW8fz5hy2mTPiRMqxkkCJF4n
fRZq4fljqEkzDee9nLi6kIKCGAV0WzjKw3/Vq1qR8VT454dsADxpImKDYMQVedIFvZLPWnGjcfg7
8SdVnLUeqBeQ8uEmdmRC5C+3Mij0XxOsVWficwvxxFMTwnylG6Xm02vzRo2ifMYBEp2rzMzgEuOK
9CEyNeBnqG7C0gCeGx3u4bZ7fxihQZSLPB3iLPXvfChPQOu5q2O5hjmKeZYX5e/xwT7qRYCAP+3k
KvOXxlM6v+T83oMU9GBzoi5RJ7HiFQJz5Q9/Vf3feR1aOmZzWUcUgQ8rvGClZlnzlAM225KhPzyh
8x62/xQ6bDwkREBvwsIh3NKISUVep3Sqir86ylsf/VIBXp4xqhIQn/h/P31F3I0o7j70yZOUqlHV
h1F2o0iqIUL9FjLWJZzfcvWLYWpA+FunXm9wchqyrrcpzSueu4AdglHdOOWYRLc6/iHIBBu24fWV
IzR1VK6/RgkUH+8yCBkQMEVn5LZpe8EP/mo4q8tbBtN/N/pmcZlBhN+WbxWB6h5u+xBzhn1la9D+
VlaYx9VyBSisVh/9x7DUlmmdOp9awjfyySjBfgK8sQ5D4xHkzl/wxzG4TbBd769SFJK50XMPd5bO
pFbnzRsyqiyoa6vEQ71vVDpbbcgDTxPrNQpGOec1XlqtZmFNWIMhbseaoZJ+1R2SXqijjSJpw0m/
T+gRQawzLg27L/I2rk4BQHuJdu5mp/WJAUAxCGpITg0411fRKT+DIUN6m/o+eO93XVeiDq6kL1Qh
DMcq3gPsUo4AZIh77EpNb6vidVbo3mF9NpwHrATkdSl6gnkjqqLDAlk+T8LsWAhDhZrMRj4xNdmL
WjrKm+RJm+mnFp4gJwuo8CzfI2cuJpHvI+V3X29M5wxZShXqGxOAu/1Zol2zff3J8nNcz4Yzuj2L
wf8idK1hxpi9/TvANknaLJUSpWzRHOmY9Z5IkLGURkYS1lxEUHTRPEdQyDOuDLcF3rACJ5B9y8B+
yJwtByB4kbc6oKC4lEmKUc0SRygvNfmGvJ1TxsiIyCfLU2zJgND0lJNF/4tvAVE+jnCLlxZzCHzo
5JEjYzFV/l1ldADyl5MJVeFCjG4tg4S0bHbvF/6eFO0NcHT0WRlPi1ACnsHh5GS0s4Sz/wIc2G92
ypkxStnJuuexJB4RI4SDR2M1L8ZrqahLzwElitNSAo8paY5Q6hsXfssLWL5YEtVk8tpMjyVY60tw
sf8p0BF+4l7ZJHcLBIT++rSgn9a+Tpy5WCgMYvENJoxcX4HIymPdeA3LUF0IdFyDT56goWChClIs
omLmhQLgsoYvi9aq2Ih16Yvl9x2Uy7FUy3/BKQ5IPsTwmurH1yvmy69SKtUwt1AVqN3e88QHqUJr
2uRFbsLfw5akzsdkl+JLL7WVRsCaanVuRjbvzecdUXxHAF0MuWC/8VIYyQaz5d6quEsPaQp4UASF
0f56VKTUJGEpiYa2riTQJCsuT4+wSfgbLggiY2xyhgYLhHx+p9pSA1PX35vjx1ju521xlU4SjH7d
QT6rRdgZyNdqXhahEoeL2TZzrecs7heCE9Da1uo1B7glMg4ZJpoBO8rH48FrDrZZuuIecuRm3HrV
E1kTpuYrVqAX//LhtvyLQGp0gR3jfaSUtrB7Smkqg8uqF/ZrN6KA8y6dJ4P58LInCwArO8YifM9u
AQecfqUSsCVUxu74KEY1eCENOk+V5430+oYMkoSy5hMDS34wIOmdywtRkGFebXP7GqakI56/WL4B
wzdBwm1vdZv3XEdVU4xx6smVMndEbKuNt3nbyy9PPPbqN9n8MzbNaVPfTyFE+N1a2wtrgAdGdnZB
FNInBHKfzqdQw2YWaa4V05BUU86v3ttIHDfhuDagpAp2agGxNM4z5cvtQ54YNgClx4MTa/07CfXz
sdO6fCu6qrbZ1Eu19+430bYSYUNSdKUu+XS6Z5dF6fp05LwVsCVifX0EkUQkQwjQwMizPalXZWzJ
DupmE1FB+Dlh68t/wmdBIH2z6n9QXwQteao/yxnBiOf71EsmTIiOPCN4NC8viOkP4YFEor6mcSDY
I/OT9XE+qCGGF0ekx17P8eflo3hShk46gCAGc7djVLz853VhVx7+41QAG3iBV7ZpxxWuLby7sSLj
bVyMizWThCOhvus67GJxV3iTTqgY9r0eOjZjiwo5Re5Nly3ng8+IuJO5tGVaUbBKDvFMtvPmxHdd
k6J2jQhQp15kbfOtOh6wRqCJq3HkyGvZgFFdUGtzHD9QkrxebD1SV8vs/RbIM5ZKLoJUMlyd0Sdq
9HnZv91o/AtMi867qnLmnK9LldjcQeL7hts04MjOMR9bwjfUtg6PXKCSOJ05RuxyISeerpsGhgkd
PuAXX6yb8fYVSbNoojFYxeQ2OusmlVI9U5niOdnOg3MB4KMrOWTAUAGotZX8VTyjELBunCkayV0j
SRn7dLinz3kYgHdUYxnkyDpPpBZHqU5vid9w2zMNXTuf3wiwZMl9jlg2G86Zn14n7B2DRYQMAkGL
pqh1x73p6NpqyMCRpCQwRSDsSQYkPs1c1WeWhjD5ZtutW6qdtuUnpHATyxmgtYlvjkkk56D2QzC4
Jb7+ItMQLOhGP1OwmZpjwCWDRQrwkxRQDkDUyapbKo5Nt5AkZn+JAwoHVXeuPtYLfQSHJ1qPInX+
xTikob8YrMofCAFDvGwQTIhIX2VZvIrXhPvlXuP7IJf9XflLGO8G5hozrXUCN4vgLkPNC8luxsE7
le9LYcNqHJJdef2MHTEne0cfP21UkttZtXFebPbS9WNDZHF7XmcsvaRcdyWgRDugvruBTCAV7342
850Td2I9dUyGznIj2kFlhuNYwQa+HZ/swqVeBJssIfmNqMRXtERVHpS9/MJ1u15ZCJsADnNiGAGg
WopSd99/9kb1ahAi5cVipr6Vs5tlswF+MI+urZjkxlD8tcydO5rg30i8QeXwBta8bqP2Fgxypyi/
S4XRpht73xOWcBo7juJLiMQS/4mDFhUj6dyq/7CoX5oaH7KflwhIAla2I0KoqEDbyMwqO4EBank2
VtiLk436ZBfeKmNP9c1+WCagyYkXG9Fzfhmz0Mw6viiZeivtsXiB+RfZW6DDugvASnd4UQcq60FN
PdayNvQa5oV6RxxcR55+5iRORDSQGzVvAc3+S72G2/mJ0wSJyL+sefCghw5SO00RmgDqDdYXUmvU
y/W0r5blxCE6wHLZsDS+gUIlhPcQ07HupO4PpW+zFSp7AWZRiiP99nv9F1oqVNddaO2eplAYqIN3
M2Ng49NZXpmNRdbd4+Z5X9puKWrrwbU7ZMQfJBGAT85ZLTwBQ+auTvSKvvJ+ixl3LxR8NDIq0QuD
pmoXbxCsQKubrxvWAHvfvNus8UK0H713zTkgzoUbBcnZeAnlnJN2kilqwk5175LRSdHtS1VGx170
NEFMhuQ+gIxo+G/ceoIBOk3hBq/zFQZBhKfFkrQCFzEW+1rhsW+nUHUW2BeevuSqlfogguq0gG7k
JIDVCERzT5jUQoB4rVXuMXOtxmqoFAw5Lvgnf8iQTOqPkNF5yitd+rpKTOzsiq0nlViHIyiJAdQa
teLWbOJ3YO6sA0kbh+1XVX0M+1LdryhAV2ug4USc8O8qa8Pi42htHFPcZgnZACDBtjLHoGj1VBqf
9qPgJA2xkkjzy8D4CaDlv4bWdV+9tIskJ+yNDzO6+0kXN5YEa7zPXOwqzPPl2zavo2MjLMPoquZL
wtwJN/YHrXXt/g8KOx8Q7PHjOD/haSrgC5R6RF5iNHSeGuWb83gMsLaC48rZLf7aBJ0ZlsW+vLwz
Gaw9ku7WCsMIDCRUDtlCe/v8OttLqvN26zPi39FyErkK4A4x1SiEZdId3SL/pwlqfmJQwNDYCNwj
qBCSgcpPgJUqiFem5HWJtPTh7CT4EbADnebwU6TGjyRWExq7l1oVcQ01PRjOcxgDXOZ+/ty0Rjyw
wR44jEuotb42wB7poXAiE+hyKiyCHZf1vT2JFWZZv1mXfu0dc0QSlOmxkwIJ3qFhH15cYGDUrwS5
UNQe3n9UEy22r/gpSNimwuUU2z4GAnNtDfD+j3EXoQZw7MHoS9MOQEwdGx/6OMFpiZ2GYGw7X8Hl
KbXoBs9eyfdb67fSbMt91GtEH48ttvW+E7qjguVzW1XjVlBsm6om8nmFoAdpPDJr4JH5oenDEl0E
0VBJiBOdAsCfFI7EUCIhDXN5RfASrMaUeuE3F0N8mlj4D6FBy2VEOdD8xcKB7pKYva0a4eBMblLE
nUuBNQooaWkTl6GgmPs9FCnGYmJV3+soCdpJmtFjYGBZxObcSn1YhW9EeAJtNaVdyvKTgNLsayFW
uqlJBArls06Rxih/XpnUzyYziknGHczYM9OD9I/PXeERK4Mh5qxHzo82S9sT9ezWuvDP7oZ2D9/a
fPeS59FIkiq6KKNILTAYieyjqwgL2dQHtAYaOXtJmIF7NtagwfPztJ591uag5RAL5fb5fFB11wQZ
3T5G7QQH6ek9qruTrv7OYhCSgAFqR2QjkQVBN4ZZu4eBnG3/3C/aF6n4BIqFfLD37Kix+ltfZDje
7fzp5YaKG3LF7ngJK/sxAVyFndTtp2WbrUCB6i4RljilnIQ+HlMUQ7B/XQf+lbhC8b01nGAuIUdX
rjgbxpfIQomRFwqP46aPanQqCsE0N1gF4UY8T1CJcsxDy27C0mG5idi4PXcYxf5PckLoy6XbOn7l
iDfLghC3xw6pFpmxRQixgot1GLNbuQrTexQ2JfIuYu/mtcbuBOWiD0lJ3CUZXmeVL2xlJEzelHqA
3sgrYEvSnP2XHvk96JSp0IPQn0isQE1EOaKjFOoaETW+/XfCfNb2jaWPLIbsnGHLZPGVHBsnngji
5iLFScqSI3/Nxie+pgblcxScqEh/GmrDFeXuT/BShek3Xf1Iam1FFx2osnzYx+U7082Pvw+lrsLv
4GJE0k5BmhIfemxmR2MOGV+Z5LIcFuvTCZYJY/CvPe5HFvtEIi47ThtqpR/FemmFpLtRBdX6e/JF
wwtNXujf7CgixWzO50t8g8z78L3n8nKfRnmAP+Y2BFMvlI/zuVXzHWwzJS4VnaO0T4oZWAJFFKpA
rcBAESriDFfXkZ5zB9gjn7A7QS4Cgr0oHAeOzQ56nlKk/71+czYHC7XvGKSAh9YE9Z8ILF/7MCMO
5ie04w8nBey5kTAs6H+VgTs1hpkRFbTVSB0d12H3ZgVIHGcx9GWfvRujmWIayoAgptymZDP8aOKr
DWH+msYJsHIk1kf1ckoHwHls29qCUQ6qz0/uHe42DundthPmI+5vtcnuw6cH8CWBb2Dt8OuLj2DK
csLKdKwrDhNw95KS0lzWPSmE+H1e+oENIpsbETehRB43XyDkV1V62iqtGpOAVLj1sNMIcIUaAbF9
GulmD+RawjSqy4syX9UAOdvmT5RYqdezo5r4AMqmPZRuRhytnzY5hvwqCJg2smc4UGbtwHhBSvTv
x/ZSAvCs8HArHkbfWf+hOmuUqRk/8GPhLgE5pOQfND9ITzfUkutiey2B1EtcoRw0+DpAlHWA08Ns
V7/FDvgRy8s9Y+HrLTPx6uJG1ke9ix54Ef2yFOro6CwoEP+lFWmsOFGvZS5shEVQZcK3c+DgOth0
ojwGikA+KmuQUxQbae/ROd5JDsah87+bxeEik1zmkGIcAVnsKVzwBBSdxkea6QdR+KPNbr4NrhFq
45xfw/U7wB066A1cK/Vmy3hIYqPK7K8GTiybOfkQUzyNjP4zuIxfd5HjyxTOSuyKNkDcUVUPw14b
z9Mt7shCtptrvbMktQ7GavyVVImYtzylb066UnoD1J5uXhqt3ArkopCg93pC226hIaQXPmrw/jkn
Cv9bX1kH6lU5HoEI5iG2TRIcUVCVipcpGuFS9YJzWz3id+kBjFTZFjgx1NbGWiKKAFl4QG1cYkVv
H0Rsd2nD+k11cP9ASyQJG4jgJBDB/Fp5UnlmEHD74XrC8X0ATDX/M1TKBsKYem8IfYuZ29Z9PfgK
QhXzFtUXKqcbRPvJ+Q97XGPrHpr+HNOPEGBRSsMuDEWudfo3tB4LtaQWw0wq4i+ql2PYhos7rkrL
PRkXdS8FETUcfMT/Pq04FGcjUuRIzSUEXTSmVkzZ2h5/cmwjkMkx8Chd4cnx61nlOPHhoHh9fUsZ
F4iUa0g4qJfscI1Y0SzdRxkH2bQPGvxZgrodmFev6QtxJT4FOGmDMo70DFrTbQ80We2nkvkRX+92
aLl4jCIu7RkH6T996nScBZmD3LI7lo+7dCO1uXsaIio9Axdu34C5nO2iTwEMGfXqXAKtQncPuHBO
GRGTgAdV2k/Xkg9CuZQeNU4eLU++TrJrEMWmr1c+g3W4mhViT3jBT51w55FdTlzYRC7Wz1aHRz6/
T8LYVW9wACKdGICNcOG3ylubeuYqtYbPjEJPdQPbV0HrRHBWLn4uZxjxB6lFr1o4t7aq7WxmXak4
kjFX3fiyDEO+AY2AJY2cLqxdwYIKZkS30s8U0AcqS+q9IIX+6/SSI1kTfagDD70xBV4M6kefnv0d
1hSucHseMSqnLd+vM9Jc6xaL2Y2Dx2RQXj5BNF/FPnrt2rv4HPcunmi6Y2bqTvMFJEP5Dar1ZV+e
07njTakXcxTakIw8hIoGvXCJB2OPJaA3oYBcxVuTI+OBZZuBAGcBm6y7ojy8lIZ10RtPVAlhIKJH
VgoxKyKqeoho8saQknCgfxfkkoNfEuX0Y3bS9aJlfByLXhpJwz6bLsjwjSUNcwC67rzekd55W4Sv
fixHFSfd6TLYYMpUr0etTm+3azc4cO00Sb+CUA1iu6osh3DwCkHG6fbGbyaU8ufsjMQipQFmYmgN
DWvIPHhqYntsy+RqR3d66vmew65wG8q7Y8vbgY5/XESp45pmmTJDY8qszcznB46mRaDIe6gUYiJ6
bP67ffzR1QcKtYMC1tzPb9UJPXyzHrzagoAYbkG0GCBQWvjpRrvNnkXC0JWEByDvrTOwWtw8+NX5
c5CK8szNWAyOBb/ObenFlGM1uLa0mfB+vXt4iyhKZKOVOtzkOu78oIXK4qO4HhQjjbkG+hkxyuAT
kjl8+dWNwvJuVVckBQKlOP2fF7xpEVYnN+wtoTvaj7vKQmk8lB1Zk7Js9/RtzP96HNHutaUsAPUY
vz+INs/DoL/3xFnZmx/cyvzEWNm13zcmh0+MD51OhStcPcJ3dZkMBjONv38BlfF0iqVal/1kV7bF
qHo1qv3S9Ouqz6PRNVthO++yIGQ+RJTihY7TlGObBn2xRCDuBiYhFMcCX0zrntFli9RPXUBfqFCc
9CAtyM1ntCV97eQnfuuKmlF08pWh0luLATX4qjfw1ukOfU0AY6xXMWLvTvSDY0HgbT6d+hhXl2JU
aa8xtmpkF/GWIQy0ypW2RCB4WnIldYkOlyOzCDgAW/3VOs796zojKscGFcBw+7+QBNfuXPSp2F81
mqD9/Vc186UqLY6HI5zi72XhlygrsOZQrz/N0KVpRqsZObYLrj6DAcbnoHIbzYPvBgVri8eBP85Q
oNUcU78VLMUZDos1ypj5315/lyapKzfhkxhMy7scrQGRpiyxvihO4lr+o+7FP7WhBlvJTqnItbOz
PYS6IEVFk02WXi+TpcG/SBrR8H9gSH8Y3XTacsQjZEh03AOy2WL0XpMwDy8Hu5UogqFhYpGUGYwt
umwxmaLcdlZnT8fIt7phOre6aAQtNcmhuf/9h4pmKivh56IY5XlVL3SqBE5ibt+zdXCEKvJAbrQv
vQq5/X6wbjZ8zJUiMnnZnRphPr+ikMLNhnDocgwymjUhu5bhAd4ye10dRLunFxqxqMOCZVUAog0J
ATpDnyOmpsbqawD/IwWOqDStkep3J0XszFmc8qW6yZH2XLjCqP/XXotreOYs3hD00IcmKwLYwmoL
d/nPzLH5WaA7zFRaltQeb+jn/Yx07LKCsjaXPYHV9b2ooBIfsq5BKYmCYXezYmmrbGRB1PzA2pUk
0pciT/htdlK3MECLpE+iaN3csSnzpgKz3erYAF4Z9zyoPNzzhaY0wbShsULIWI8XWNTD1yf1LfWh
aqUxpUABfAUl9vTgI05V3GEymIfyPRxJUzY3iEcMelahEq360TPt689GeYan3BdV3mlGJNzOH2ZH
6INbyEUOcsjEMAGinXuTXigmTWneB+l1x/GPpEJQ/o2zY0znef37+TklC39v8ojGbW/HO9D5q9KP
rC1BVU8U0mdtRxRfbOUoDby9LYn7R81oulLU+5GBoNuIPS0eaQATsi/33RGI+e6JeduoKDZ5gOps
Vzvj1H0k+zUE5I53F69aX29CbQ5dsuL1ZvA1x4R/vTJcA3IktBU7Dw2GMtfPClpZ7qxmF6h3UyaF
9eehX7nvaCQQVzyzsGD3b7DRA1V5Cg7NSBcJIuFFq96llIJn9jn+p40YJGhJ0MVSypoJhANBc9Gy
vlGzhP5mBeDo3U7EBiXj/0Uhv4ywHlRFKP3mAOPHgnt596o2wu7YjGbmllnsl0ErIREIxd45RhP+
Q4GnanKYM4fdtNCdnHDUU8INlGHc/WdugTTcTGJWv5lM9mHOYma0xXcK2lns+mkVCB5wH9OSijqP
pQlmC8JRXeXtW1HqqCiub+YdE4wjSQfCvDW7triVJmAneM4nuPC57mfKKWE3BzLJWjBDwmJ93zJm
pWhCbqwis8xq75tPQ86TrVXHR4p0jjXDAccMYjfHGX8PY+nfox1AJFgPSVJm6oUxaeJ5ouyMKytI
/WsztIi9661ZriyNakgaQtqRCPz3s+XAiidIzhgL/y5anpaADAazDiTRZEjXosKUyGycoP6SPd02
Gf7re7K03e/oP28s2tjPge1crocpAL2rCHwgosuY7UQetUj1s07rPrzM+5yPSl2A0U7pbbnFV+Se
yAgWPi1AKEUqSj2DX3lBj8/PdxSXerBmJY1FLmlFzPZaH+xTzie2Qs+IU+qbEcuxpD4vYRzVtO+8
XOlfpinPl3OymLT7zXxIetMGeRxr8LayMRt208kz9h6AHOHkD5KKq5JkSVAsd1O1wsZTS/BsOcHs
y9wCwzccU8yZleQ8seu9xXEQQMVtW6tRK52yL7qb8GhhaadvJhiVX9lNJosVBZQKycvjGYyxEQH1
ybe17OWyAAOEWRB6dGw9jqIbeoXQo505IT3guEpR8QKeBh/bwydtKVoxXtw6lHJVCnIBd0c2CCVE
SoENY9OXwnHRt82l41iC0nNCv7EZ2hfywSly3xAh+psKVSIGuEsRvTZsa/yvk6XcKnBR9iGX/YlN
18JlQh1+y1035s9ikx/fofZXmlBRP4C6y/ZOxjG4UvhdnSrk0vwiqBCabxtQuYvyOZfsJXOjGydr
MDVJhxeKIYeco9C1VXE03FLa1ttPpXhssHL2wZH7ecNajSKcQjyT1CR1OakmfmbfeHSA5jxrmE37
xsvOXqrmMJldkJg1RqK31zmZYT8FnbSpIp++IVg2wg2yl9NysQ0fcwQW+SUfMX8KklVyzItQuQcc
McAIMLexoDX6tEX3cY1esF4ChmKn1BwFZ+RmB+D9z+LpVJP7Ar4QERSFBc2rn2Rs8ggL2a0R6Ok/
DLsi/bjJBS56c03jftdBLYawLNGDQO5er1pJDtxysYZCvmz34gu0OLmD4313MbtOO8CjyPn9iCUJ
i5ENfj2Myx1POFLJMGZS6tAY0LvGMu0I8flT5smX/M1co12QT4Hbuu2wScYP+p4wh7fD9f/gC1Qi
Y/64J9t7WE+W7ax0epH/O3Ek0/jTr1BWr+wRIBSF5FFT420we5AX1czC0V3X9Bz5MagcKXf3j2sG
kbiYdik4w+P6g+qsva2BfxCUhITWA9sakhTjf5qdXXchSCOiyvzTVkdQPiCtcQY+3b0TgAjikNNm
SpSdVOXYIayixwgGyyRnT3rz7Kdhy1m0OrtSNtobYdbCfyc7avz7rc7YSdIo43k6JGqnluETLHAk
gRtUlm1L53mx0M9h52ZBwLayWXWRI3DeDsAHPEmHYmR1kaTDHbSoaI7Pdrg2JdwcTOWzPwF1qgKa
utueaVibmsN6pn0zpMvFq31bBwhUNO1f/TjKGj8Gw0FKCHYjCbGNJKrLVcd31GnhixMvfDcEHM/m
WAn6QXxlcUBW5f9Bh0rB8jpr0EaHKoW3/JKwMWEmleWBiEdnOfPMSlhFqS9olMRMDcroVzds4MzL
CD31MC5Sam7gZWYKn9+ROqBq/X6lyrjMTWohzuF1T0s2pg6eWdR1j/0/jAM430VgWqRzJbn85+6H
QYpYSexu6hfIgyOa/o6HiR8XP1FG9EvGnfCMVMxDYsQd5CTDBsjcfqZJimwXTKbzo/dKw+k+4o3N
erm1Tex5GUxYzC/SXkXIZtF+/NfHObjAqdNf1AhWtywkppIggeD71stvfyuPaloVbbnO2lPzcSlU
AksMlecUrEXAhh9ddBicP/yGjGW0hBOIYO0b5GmDneZCkaWblusQ0VeB6XY9aqfjIs//EGr8SVYW
GSSB/tR2UVoXvIE3VYPqmB5qwTgmNbkgdoieKjgjgNHtvhxnHH872ozXfUyK4gZ82p2jQ9ybCQbT
f4I4I1IjACBl61tZRaWHq+tC19Uhi6JXOzZQGX01cP6ldqOS9c6tMTOM80I9Uv/TITnN2k0cPdT6
Z8MY1L91PVj9av/RWzNlHDWhdntac0Azg/CV3mqJOibc8QXq1GH9hPKp0RFx/ikt/EMWhtpxTmHu
82h8oegG7A75Nv1mXhYnnIwkMuIjsF3eO3ic8TzUsx/RgErWdAwjei2oHOM8ocyeVPYVVFfj6wPw
rAY/whlWcknQ1U6giSMuQbLiOv0bTUNOFwFg0uaHrSsVlr1csQVw3NCBuyxslcjp6Xzzb8GvZM7t
X3S6lR1+JSqW4gpFjMWo/LVz6AHtTd9EcECjFIxFtYUGohzuyhqvpPYfcDx1dT/fUYMOOEGJmhCY
keZ/uWtW/VdFKRPafcR/8poMKmnj+d3QfUYKkG+y3HKAm05qsiIXjx3Rfkfes2WkpIyG+PfeZ+3b
Asrjja1Ipj6h7tNGj3Dmao5LjJ2FlbmUisMzwUDPuUWa2LRwrqjZvAjAQDdisqVyqVM6YbaHBBqP
LiXNgS1LNpR+m4VzHI8wA34DJDCFjqZvuzrhlsTVNzXHW0HJA435Tb0dHKsQNiLew9FEKT6P84ce
ZN/pqZVtQfJN9w0VPCoJwi4pePCuDCbCtrCLsG1NPgYcb26C0DF2mJC5DkjXSeslHapflG+YkZM7
84EcTdaKQoMY1SGdLBxjvOlhVlsEUaRFR5CQKo4clSUDZxGi/fkV5lAvfVW5mMM3lREpyN7u78qb
pszfLoAQg8mhaN1EYbwGQ6ZJgxVFax/NXyDjgpmyYU9pEwVFbKRiYVP2eFEPz/vpkIPR02zwzDh7
OgirTc/lkXCq3Oou1atZnAv1LXZEomtFhhq6TY9I5cA5zEsd8esM9hrXHY8E7Ax31vvu9hJADfpx
y/cI8i6+KtnRIflXTpjxT3U6zfLEWtdN5YasoAtdplFOQw1h9g74v18kYRz+PwTZD1GqzYwapAxe
yzh3RuCI1ABDZcBCVLKAhYXJpRgboDFzUWzlWbfCZJBtdqeNFY6qmoIfZMVebSLoxzDyWKRE8BCC
bzCJXagc0+iQNUjosrUVTsZv/eJ/XJTm7NFlcpY7+8hwc0ZUe7tChUsGwqcD1aO5vsP2kpBqRA02
qLPUT7Ovgox4hStIrAG7Ihz3WMQaibxwqcKSbcvBXMg9ilxZHHnkypMlGbffVE7Jtrxobuf3wxQl
p2M0MJ7NqpDA9QYD0p4oZMvf/l+dwtVPgNKmYHE39G2LgEsEyyCroPH462kOBbT19cujHavhvRKa
uAVTJFLULqwGjBG+gxxtgcEQaXiME/U3Ll3MMC4W1RDF5CG7FoNTP5j5T1eX0CIcdWmA5ovVlQ43
P/1Dx2lezTe6lGnnKT6o2cWC/uqtr2g0inGx+EfzfJsgd93hQn3h3OvPjWaHve3vYv3IW4DF2TjH
s+aHaBHByYtPe3DmYrAACivGTNiCiuj5oSql9PCZx2tkpch4ISqlXvc5p9GO0SfCznwwyWAA7J2s
E2J++b6Pq4TrQgyLzALiJsPBwjlhaRBmuitZNJ1m2pv/6bdfHfKN911rHkMC//HJPkTBSDxyUYde
1WAlUtQ1nG4T5GdDQnSJ1zYzesqXaWvrmi4fpuSNy4pKsYr+XsoIqPkeSYBlPsDn8Tk7UdzPGFwY
7vVTHAV5H9LeQec/SFayJVXjQqjCszbzyr9kaHs5wWY9RxCai+RRYAHlabyTfHbN1FlMaIVnzaqM
MUtaOrFLD0oRhEkg9lku28hgCT4WN5h3DbY+47N8ZfmtzQSpuT427Vr+0FaffQ12Mc1j1t41QOyd
AcdG7ZugZ/TAoUZEhDrnvNahKG0S9mNRw+4O2aDbv/NMSzj4qZ7+5uIxUpnUGKTqN9xBlYqmFkPl
2DZhLCVmmTxemjdb775jUyhSxcEllrVvNE1TFHHkF2oIg6glNgT0asIi1hVqVqM82XXwsgKiNg+C
G4pGTnEd6UfPgKIluMZ+L9KcdzcQ30TYAEQi7n3gQct4J7QhipS7379MhD4yQxsb4KYzHrh8jdbL
WWayRfKk/KzVm3AojY3QmFRdb97PPgOqmenDEjwOtjlLpr1f3Cwf6T05lxiLhnI+O8l4P3Y3M9dB
jsiY5EKcQtlJFVIy7Rn9D/DawzJyH/5pBV9HwQEfvTQqJa/LqVT2mlRuKwGV5cIkn1P6mYH89Cwc
8k7xRE7RFGCH8+QrFIC6qbZZrvCoANf2DpMXxAzBBr9OQO761CHKa3Xikj7pSER49XI0JtIbxej2
3DXSh7/mhAQ9H6aHEDOOpsgXjW9q8HLn8eZZaCp0KT7oYjywJ8QtvIsixK3HIgY6RfbbSUXrg4cz
vVcLDr2SJ0MWADYS0z4jlx4NgAOGtVokfR1V5Cj5tGATNrn65tQSlASaAEltbmDQE4Leth0DHZy9
buUOUIUbdD+JBarY8f1WdSpd3V7LJfqdzeT3Qslz0DtJnEht20D4WMCt2bd9EeqExcZ0B+BS47AG
Vvh2d+ZcE5X5v351/+EPSvTYfWDV0oYUJK4Za8+bA3/cui+RsgdCJWtSu8y3lNWrQjbqUIp4sFj7
7WPgP9lFQlBswcdK3rBmpzU3THYsnxMK8mArmLJUxYDbTzfTXO1FQCVB5ooQ4azAYDopUtay38CB
B0Wys6mh5rcE4npoM96fETd4xs1GEd3M0b5OIC9brdFgIfewbb6BR2rHXpMihShpTqJ/Ip9Urri1
CDZlRUphvw8XbIbjVJhk5YcxNfEl51PXErLPiKN80L+let+TcWspqJf8QFd3GiEvjkbbFZRs5nbL
uvk3F19K7RDEY3BQ8fKJqd9iBc7iRA0WC1saFeXzwfY+IkR+qtbdGdl9GEh49Iv9153Yn1VaiW1G
DRYghXqlAofXuzCA/dl74Mh2Z8xw4YWTzaOKefyt9UlWuemU9zOVXFh0QziwFqNIIJPUUkDXyfxi
MEqTF5SeZkHq/qvIJsVEcSK4rXVNnvNFnYsm204KkwBS/mv7GnvtyZmZov/drpJYcu0GF0EL3qhT
N08clMyMp76m376QXgmZTcyhVMk1SFcP8TpC+UdDNG+DPVbh+QHIf2miJ8N0Nwz/ZsRhYR+HGyTi
UQoyqGbB6v/5YDPpOqxGxudGg+WITzSseu5xfQEvj4tsOdVKeSDWllZvFru2pP48pA9DB0Km8fg1
/LNIfhjeVkgQCSP79kxrn/vJq/7mTDij/xGByRvxZ6N8ZDBkCNxrbNEaCYy/WShDStHyXnuxd9zn
3yaDIiHIzSwiwbBFWBDGVCNYDYy13sU7A95xbWEh2WK4/oeOPKKz0/VT/TMdM0C/6C/utpFoJ3Ai
wEoTdW6+FwgTwUyfJ2l2anOXKIOdtg+CS3OnWDDppl0ZQi4nxYGzTSE5ymUH049bVX8noDWeQFVk
5Hb8uwlBgkNctevYi0bzOs5mrMm/imdiQuUmGIihxbB6z836BOf+WtMDucQvDBOp9G4ktV4lWTy2
mCfI1t7lC8s95v3GjIo+GAQ3m/Nc/aLoKGoddFofm0B76EidW+mFXRH9Kv7wLiTWgjUJ3hYjdpD3
YZqLhyKPk0SdyjEHife9Ph8u9y3/vhstt7NpziUBRbUaH5vyHqyKQJhv6mZdm24aVY4Of9sGkncX
7EK1aQkDsP7qAZbP4bIMsjeHSU4ZvqXebRNxyLGVD+/GgNQzbvs6IlAr8QzK+1FkQLgDlbph2Rv6
wTvuK0eHbiGDvxexfxKaQM6mpJsTEpyNPPMVU0uUMF24km7IpIH+wYH0/nSX02mp5cemcdabDTEw
05sIJySasWEbWZgpf8YqY4+pamkvH05H7JYs6QefpddYmN8anrbzkm5AYZFERqZEMmtfzg/QzW31
ER3D4hctysX2v1OoXp09Bw1c9JvwUzBts7xEAUwuwWwouKBDmGdKHN6JDv4MReR7bIGxZWy1e7ns
6e6DyPL9gTYf5T4vJJ7I8vuN5Az2NDSz99ZPbbvjwnUTxNccnmE6krb5GAlTBKqVJiFJ6KsH9sqN
CboDmqU/buw5qLkazfNJyP7xUY/D0cYURSUeZwCFRvnQS4CHpoy/xVoCrNu6bFPmC1Y1emoQPEEO
KVFBQceEgPFVj8ZrLvNRuZP5e1DfN3wMQ8/MiC3gPu626NKO8E2xt5DPrgkP2aBbaojwbdlMKK21
GmgO4ktArv5qzoAMDA79Je53QvqknKE25gF5yOdvU+pFtqKkVBmboaaSisF5Fp3j/WD8qu1A6BK6
zwOeJY8DPapNVs3IJqKYbppXqomxhd4mJc7jTWcfD0MauGktm0mU9z3t7YrtIBOqc3+4wYp4fmwy
qqzOURcC21v0PaslZyvIg+OCnTVczWC6ApeM5Dgtj59vlSdy8HIBDYbDXM9Qxxd569KpnICq8vG0
cs1URWjuNEUuKC8PS3GXDhiE0Rh2D9bj58/JNLYN9WzHud3VrhsaGmdsZUMSw8Qrz7XG2F5sxP6W
FxdK49RINzcgO48o1FuYMV1Ib3HHtkApK7rJ1cvgc9NBC2Boe5ovslnGHYw/L/LVujnIlHh/iq0N
/Dok+uKWbrBkA4nBq89ORyWPJD2rGgG7peNSN7qFyXAiV6rZN3HWDG9Jq29dgVbLYlsU/wfjL38y
55Swrl9yrL4MSOtTec2KtE6B9p0NEtoZnppYeT4ey8zcE+DGmXFAjfLTVPlyz6cKZOPLxGDlHK6j
AIW9H0TwPmB9mUeiEHc8h8IWLhqL/9vFNNGaWRilNTKv6ugVlczBCrx/N6EtHh0CevTYsKvuBnuI
IyBQKpzVImQTLsU90c8g5JC/9sETHrdRBLTEGjo2FHZeOFE/DfWeGWYs9g41pji6xskXZ8063/y5
+9kGld6iBxzC0JaDc4bCJ+WB343f2ko9n7TBD8w4T7ce/X7kpmo7LN6ASb6mBuA4vXWEW9+7yLTX
pYRkPHw574B/xe00KZ/SW5FZog1pBnNJrC1DdS8QXjqJyxvGJPBT2m52oad4E3MSAh7F5zjS2vmF
Lj58p0eiHPtON80N6AUvMWmuPd9fkl1pTikqLTD9iMVSdvVCD2SqxmiCoaBZyoTZlT38jEeA3ozH
3Vhd/0aw6ymwO18KQzN9VKCWno2Ihq8Ti9erLaNnmGn38hwpk+Vhwcb6Ih++oyPbI/Hg2rrdgzYr
KHedWZ1aZPTzm1eHI349h4nkqWaMTrC2hyLYAL90vqKHA2fXUU+rGmXISSkjkcFPJ6qAb2a1fjm0
A6eKHwEk9SzgMJDyfgFcHlz1r75+Pdfq8WYmeAMzI1NwdACcVwGL6SvYEavVT8V1C/Obu6G58gDB
XqTisMZoHwY54XXFDuCpJk2OEfjM3F8cwlCRjDFiuCpF51gI9f0mcuZI+5L5uEarIhPitonVTStn
AhCUNW3yIW4hyRmF21IflCS1DrDTEhbxYtZ7dcjQ0JDwDVMhuk245qellJ7zdK+dVgJYWdfza0kE
fm1EnQDD+3vKVjXKiCaKqzzO4scIqxIYHN3g8DyYzfL+f5xV9bMUruNDgRmnhEipaY6tl3FfrTZy
vIv0wClv9tiZlaDgvDeZstz6xjbxuQ7PiK6mKVegK9VMIVmvV8rRNgUDoXSQ3eor0Jt7wY9fdQCi
3F8OljDPKLPehtr9vM0DsfoD6fZvEuMeDd/axIONGzjK3dy0R4qGQtNYjsrPIF6hd6UFFWYmq2H8
Jdcr5VAGKV7tclc0PwH8GNFx2OI96tyge+lLUi5Q4I1N5KPE4cmifxfBDtk/JFkSgPdxzywpJLK+
9cBaY3S+3UWM3U3gf7qmgCkr5fBVkwcdbpMZjokOuFu95zgz5AD9HiQF/RBrwuKDvfJT9KsW/P92
IRkI6DPkpOq0MLqA4T9kXx7lRUds+djpq9/OxKU08WI0Z3H7tKqZAlFXEVvykHbqWL04uZu/MZDj
3HX38/QJjgMVq5om9tDhaotWsHZ7IvFPvI69CfSdoLsYPtpbP/RaZUOGkQ5itB16SZLZaiA7I7xp
dodi4pciqBn+EWmDXFgAaAFLa1fX+/tDR6R7yGxraRTt+hYrRDgdu1cRR2TKAnqubRnZLst4qhgs
jNy2k7+9UdJ0B9cB2AWLw0KeanMh6hsTNVA46oJVJWb6IPr+u1i/Cg2R8ARr2nAICr5oarGW+bN8
mfMThd6acSPnHPUySVuxHsrXC4EZSW1gdfgv274IIgUwVueldukcRtxIPIsdMJ5OhjfEvw+nduvh
BVPMMUe9XOnxo2YJGquuwrb2NYHXeGHxgltLtyQJQZMat1IOdUrIuyXfpPWteol4ZD9gGmzEhDjD
9QvZBa6Y4auhrRXde/uxKaqwJhNosn2XwBUUXCSE/p4Le0p0gp9/tgDHFxRn9d9cTO9okJqHBLq/
JpxqSs6zs6lbj/v29Y9LdvTdu6Gmju5GBU8kKT1fecDfuQx83Up8JMCHSp7+6ZY5xwvt1FDSgHGy
6OYtNEggAULAlEoMBaqr/APCAgsYGr4xjsqVLeRKmhbV5M524690Hup1d9m/OXqD+WIWqHpdpv0r
mBbYHlUcRwQz4knZrBF3aY+NiD8iMfiIJVL6FDjx//ac/JkF86WBfCRuYitZEJ7tFz92VGHdubfF
utx3cvuoLJrhsiSHlca1NJ3cZxKFunMr6jgn24Wx7WY6UsclpZ1068iChROOwBGMYS3e3fXC6ojX
m/m2r+diQpx/qojQOXvXqIVAB3vzJPrPiCHPWR+PrRkhRzZO2HYKq1Lcs6iEMIu/itw4I27U62Vo
8FzI349C8H5yPcVeM9lfDy3j88qh6spQ8D/iq7BlQSt+xKAp1jdg2kE8W3unc1POGy4wW/4ZFQuA
wb4ra4cGd1K4/vzTN0KC1sgavqx2yQSaMeZOZvJgeCw1xtEOJ8zfwmx1uDw5K4W7q3dR+q8vndLg
71sDtMHmY/017iKjAn0upbCLTiYNnqoYx8DA4/Ds3h/5jS1KPMqD0Sibx1LmJCRBMZY+AFkoXlca
+qgppGDKdhr5eVe5/kfR/zJzfdYSbCFNm2BMkgxTGK75HtgcSDtdp1a3XAJubjE4RdV4RBS2f+zG
NeNil1kui5lPDgRuohPnslvB0/BBAEJ4jJpP8h5Pvpglr5fGBCCt0EsC2Eid1ifXfm0Lq3gWhp6F
BZBurWp8waCB93DUOO1hnuMGaivXpYhLnvaZXMEMElfcg467XeJRUKOLGcxN7ZE/yJdj2O9wt55s
SgSYQA2YfZdDRfzH90shBQJHEV8SMpU78+necQspcdYzwdzuQWOWSySCyaelfAnVSnVvNdFXl3OT
cfHW05S0XPaKx+3jP7szli+sX0yx5TaIi2F5GpOem8XL/2kZ332sntVlWGAc/Y+GetrQTC3cUYux
owKuNtuiITXtzw5Eh7aRoFjQH4kM298YNnPeEuN2/pLgtWOHRy0uXpN5OCAgUdMaunLtlFs8woCb
C0ciIiiuLU/SdD2eNAGeL1n/aogDu5rjP8rYqe2NZeIacr1zCtjAe3oU/kMWeiG45Z1PXftS35e7
RjGNfGcPzoCoXoU7zbxx1uvy4b+bpGU8Sz0o66IgP6d1YrxmLzYhF8UQiNuXp3GfRzv/1RadNrk4
+aW++dI6Ngq/dcQhf2Hb37WCf45iN/l1y+SiD/J+1lDmaZBXKj+yreGOhyaaLKeIm12Ict5h3Hdg
EWlC5iiVJU3xmQVdci2PBdpgbJDgOJmVQj+Td0w3pcOIwdcHsknHY+iDS28mM9WFgH4dwe+KZZgx
AH8fNE1lba4rCcohJKiuwq6C/iVz5bxSGWOpu1JXRg29uAPNSwdGdxXunN2jLOxnE8xaJzl4J5HS
Ykh36Cg6nJ7fy2ptuIwZTGHHnL2x6Ky05ZCyOkdoP8TrjJ34PsfRbnYE+8FAMYvt0s6cgxZ8aeYw
pCAWEbe3c9RKTCyKJsw1q2YQ5Kn6CDyrkD90Yca6a4LIsxlzHjLInydBEjXp2ukCfCKQSWA8tSAq
dYtR5POtxXhGxEW8oiYtrNPd8iMv33zWBp6HaHAfjnxmBbvv1vzG9u/+mVPit56xMumKL3U416lj
6PELxSY8WzOD3nZ2WxbTVTYF950gA5FtNVAu1LkU0XG2cPgWtwDNt7gAHnu3kWXWG3gexdremAzx
sG2AS0mxNe3jbtAvvuQwO2gVZxmxwbHJ7zg+nR9wcyHl2S918oDXe6h0qEDOdcaCrP1a3wmjqpcE
aKYFUsQBEZwM+DEW1USEPGoHcEddsNh2QopZ46H99zK37WQg0Bqp0LB/ljPdWGBmDE7zq0pBlQ92
OvNjyyZQzBLszdzDBfGTjMmiYy9BZ9AR7uuDWYVisl8izCnNOgnpRheOfa+v6Imy4r4BJAQx7YmS
/Qa2ZoeyCGKe30Urg0tggG0WmBIbPipOPXlgMxLjKcaGTNu3gwtGw6yLPveqfcwpvJSbedvOeTu+
lSICVS0cnneGhIliGLT2lLzNeJVt5V/iYLhlzAfPA6FgYgVuK9b0w4IPiMoQviuX54oFXVeRytoR
tMG9qM4/j440o/2TiNNTqspC+k2Wn+MM82TnD4Rfxlt20qd2qSni3D0VqFM83XS2Zrg8UWIy3wTX
DCs8c59jxjqf378w8MBDGemTebBVS6WLaOrnTuKJ9/6lXg9F/kmwNDUHA80IGcpR7Yem0z2ztZmD
hdzjI3kpBuT+5qS/XMmB81sM0g0/AELRoROM14JxTXbXyVFwrGcL5GoC2XVaFSQKP8gGzziEJ1DM
jMdjhkgiM5aivAhZyccuxzOukgLfIxyhbWv9flh1e0VERYwqvp1z6TyBPl84wAB7HLog3jMJSbtG
yyzm97o7QAd5xMh5jOYkWXGdRCv6IeyveCC7SGRQtRwhukGTiypuY9E9xbUvgBk0u6y2JqfEcUa2
3+gciXwTEXGzeJhoK9o71QXlfDQrw3/eDAbePwSIECNR1dy0atPwC//iEyKhW5ULct9YNu3OL4x/
/uFJZAjSUMQURogp4GMiU5ihUlFOtfJnXnF3cXxCA81vPpcZBLXth/8zGSzvG1yzVrOTSTga5Cq6
hPx0cCw1ipMLLR4Hu5gaLUpco7/k8ZDpAsLbmPOoD8BfU0faqoTjWuGT3jXyDcz4OYuezbmGAK56
yNQKXo4l3VhrXEnL5wk9IEw/xfs8H6FfP1soLHNJDQyfACHUUV/sxYk65zhPOUHGXUPM+DnaF7AN
Hmi+3pRzoEs5BVE53kzln9JDYF65VDC4lHNGggWGhcCl27GBy+/mSdV+xv75XaZNrzxUX4j0szcd
wii0zp0b9nPCfMkjaGBMvIx+Mmpql6H/7/iXGyrcp95/rzMo/4orKbErwsh2P84H7KbZQ8/gxvJK
Zp3XTuADdUNNAwyzfCnuQVlk530LdtY4Y7pcjTBegZhrgmsWaBOma7mDCIYF6ugHq0ZpLJNTZ0uy
L3VWssSHjvg9Bej9cBt//p4kusH4bKFLXyq/WBn1LFhmsybTodZ5KcyHWD35UQA16ApodZB419/6
T/tQvQn+lICpf3eDuDwZIrbTL79ik4wkM2S/10vF+aeC9y1WHwHmYbahwHgRW8QOzKM2svWIwuN9
TLodYrETtVLMNeuV3C5EBc7N3o8ls+/dNf/40M5yb/1TDxIIYlt9HxBnJkgYGtaXm5SWwLkgmiye
u/OD7eCZfMraF+YaoCx3+zr/T0dDPs18DHqW8BcWCYuo+rou9LovYMEnO4vwmKx0l9gLO3DGqDx8
sVb6C/1RdqD7vf3DknshVUEVp/tqGldGma5ToxujwbfLeSoRh5SszBDWQuXPfB3ROM/8gwJSMdwh
74SrCpK2m0qTTf953MqfXV+HYZ8e8oym7l3ukpLIRX0LYL5esocQ0iogSiE660d57o5Hz0qTx7mg
kNfjQx7+t1ksUb4rT/OSYWqW8TcaryW4ikKSQ/rw0+2/nBbCWZNKvznNgGZnotggIXDnueFC03km
JTT5QrRWVPYYLkwgdu6c7ntyUlmkjI9io/h+jAMzggFygDnnar9ENJzYwKXvgiWe+IAkqobMvdYH
MimLKdsSW0rcwkPlc1pl/W3+vWLQPLABkPjBs/IaCoeQz02ydsKIlU6mQYaidFSIDst+pqo7LUAK
TKS+nge7ixm0Wi/zroefLuVFPTQ08wWnkZa8TcI41HOsMUmWKVi7d8UhwVRAh/MlAlTjUcyLIsWS
F6+4oGcQFqfSfUNBaND53HxK7UdunHc5Qyu6TlNxHa0lhHHfdf0AfC3TRHWSrUgpiVMSqrnulpy0
fCu/9gJ9oVHiLi3lYc/SzvQ/vdb31qUO/ZE6AbVSsIgz8SaSYAWUgZEFt97wCawKpzRviBARbeO9
lZcKR7C+2oJtp0OTgiGL3qmZy9rMc7hlbTRydkVPyrqaCyoQTQLbP4EsbiNJF+oQd+Yv8Sqr5nDf
bM5UcV9Bw9OnI2OdB41x4PxZWcmiDO9MCX2oB6CXPiVUrTE0wE3/2XFbHWN/G2pIAfB3a1SQACyC
SWI1UwOmnNmZJgsQbSl4C12Mgn1RKEtRdmJMFh9wByst3myVdJHtZT36bTLlwiowWcHEhpsiMslb
osXbKBG8rDVAHoqIHVVI8e4Rr5m28ICmt/DWS+o92WqECRUfsX+zrMmOUlpWmvikY/426qbk2Eb0
14RUrXJlHcpwlbANj26tHrH+XwTU6Pge3UY3KlP5sSKuV4zy5PbPZAeNDHl7Gpvudx8tAp1o7W4o
TGam6y5Lo/zFx3MycPJG6SwF1cHLAP1CC/5WrG82ckTMaUb8he1piveEAhFzrlinC6eVb4hnLOCe
Brn9K+MW50tGTXP6Tt8/iymWjL7ig/4/MLOW6xPtszHGhr9Sfb83J7x7xV9ZLFNWj3EciF5q17Bf
dMZFGfcGc3Tgdz7gRO22SjAW7Tu+GMrHv/lmGlok0CZvsVPjw2z135SzH8fVdw/kyrFKtG6Qpyjk
NFxnRCpJy8rV0k1Y3tdea+O1C/a/7t6euQ6DqaHmZeyMuUxGxfwi+tOHePQg6PF9/WgSL7CjVVWU
EFa51KqVXlVZvpqy03vP9ySmMi61aomBbtx/sjHI1E89/6VOHGHj2E+lV+F+NCV4Ny8Q3NY9T97+
qpvih0QtYlDegY5014qVJahn0dvGc7DcssdvI8GC5XBX39847PfzR9berxDEalvEPwpV2F2nQmHv
pOipjt1aB8/Std60nIt+q4SYciXmSexa1++GSEuVTiwaB/sIRVmB1NSdqcnLM/nWocgCjEn/nIu+
0L5lV1v/NPv7KX4otqqy6jX3vedZFhmcSVbXtCSEhJxs5fk07G6LGJuVv4Lo/R3c7czZNKq6l3GN
rVCrmX4AZsihE5PYQbANlQ8hOb2kwSIeFaZoQ+wiQI1KQ7xMkxmUAH5K3F6mRMBJtmYFdwruudcE
fhX+8am2uz8x3SfIhbo1zcDxKbANHrIWh/HYzTmUN4b96c5EopWz2OSMSxblBXJDbQiMhCbqDWDg
5XdZ1jYr8dxSsSrBb80oSOrn6sS9RXOnev7I2pQIyByzeHGe0ElhOJD4BOJC6qY1jT/B41vlpVGw
dy0FfZWizVJ7OhsYm+H3HeOR2VLYpC73DcHwiXaD1N18qj2frvJ/HthUzLfWeRZNUViBx74zzc7o
nl2wRHK1i1EjWq8eYJyoclETKQmaGOVaMMl0l9x0ykXcBxR8E22VrAvY/68TxVhf2W6R1ldEL17J
LSdgiGLhLY1ZvYQNA2Ilv6mPVU7S9pJ2Uk+JPwXE/IqbHaLjphXcSMau7z3jWOkYUdmJE6xItEw2
Dbksupqbz5VI+l3mWMWl7WhbCxOs+WvK2s5/eXvYg6tHV94b8zsF3L32a5+50/AGrws0irDrn+Us
d2iZ5Kzhy7ituBHoB4VfnqJfDAiqyVtHL8Tfg17EgxZCKeHW/SSs801NeNMmBGjyySeEzYiSRbIB
9O3BTSbGMLRVSZNDYmm3nvVwHt834FSJ5sGdB4/7WlGgHdhDNHWfFTtRwoFgqrAazV3tM2eyvHEf
RiAnNE2H5doPJXY5TABr2x8BO8UBfs3WB/LvZrnHVWdIA42NJMmWSwqkfBGn/RrCtjCreTA4tCFV
2D0T6ERHGH4qrRums7SH5Uzu4xRk1R+QFccEoyFWvkkkMEr7IPLS6MQeAA4hkp1HlzzJ/xnKrFzk
WD+hkSwInRngLSMlZVwWlavjXqTG8n96UBYAHcJqKE+zTt+FfV6H7L0fKTpjAuhQl0tAZrMX992D
gTZzqiMz+biWWfALTZARwAK+PJ7PuELkCZ3oxWdlVg0a1ApkTJ0opYG9PSjiMpwTN3klnQ3cdsqj
9YfVaJYHxKqM4CdTQU0uIM0qN6RwECo/ziwYsbTOXt3kTpEO4nV/3Cj882fzBwrGjLn6t6zYaFwl
68IwvJJnkJd6QsNJba0CH4LWf7r0fS1FL/i2B2Kr1hOt65QzIHaQLT0SgSGYa1VKRcVYmieMAK2w
AbMl4hZ24BgQPXFDB4XFZc/PjYclaoU5dbsyEi5PnJgI8qH2b3RKBArrhj++Hqu/uKmKCukDV5wc
X+cezgpIQu8eoeC9ladPntm8wLyiosuBpjUJdk6ebu9159YCjQ7+hG3AKxD/FcVK+bvCMdAsbPAW
dpvBQIlOidgcl9Y39kyaGuHr+9F/KxN4NW6qcnJXrWa2N0FGFzVjvn5l2SzsZN7ec2rS3ZxL/Zi6
hXFywulFTTrJ0jKIrYXUhAAI4r6opWVtqM+9K9XrbkmmAReV/QSb651pG156B9/PQzzYXKqjVbK2
hyPAF1Br0O72vESZSWBXhliDaQ5dwxb2KNV3J1XCl0ib7mYhuesYUe0WwPnhrtoaY7miAj7NF/JB
1mg5aAEmb8/9/xzBL7veJ1mUWbeReorJ9Uel7mt6gavCB+QDQ7uBByU2G6iBsFhiYehpVIu5wGbb
O4XlnvF16PD1WA5BxGFwULkEZDY4oxmQBjQOdIcXR/SOSiieu5rD3Q2jHwYcOTutsay6jx5kR//u
b45NPpqLjyZG2H9qDO46Y8SNSiitPSN1GRSY/xr2ioNJk2uUxJcoEJS0NwA+EmNt+2oDNsj1X+Dq
6LmQ6Z8fFuoYq0KxP3h2CNT55g5HyTBd7b2hnK2UfasOePp9qvKOZYTgql7rjJGu6DnAUUi5uV30
WF9u9eo6atB0OsIL+MAbTF38fOiflDUtPbDuFRBfOUx3pfTD+BKgS0Fba5O4uWMNiqTroBw8r5qt
x1wb1tE7uZM9Nxx5762zshO5uniC4XVw9NvlgmLYxWZqRg5gPnc7hBW9IdHFS5cfEzZKmusFB/2N
S31+bGUYts0SB8Kz+IF9iGV9D2UWM7XvkrYmwoPJa8u1adSQPmEQvUZLUa/YcuGR9hXczC5/PAdx
kHs1S6fPfvxHk6QJnRSD6sSk6cjRKc4MFjj/Oxtq+89X4ll/M+cxXcwHISTzs9qbikk6ZQ4r1azM
x8LgNswI4jdjmPKhdVNn94WTmd7r3QrCgRfGCve+19qO7Xs2HyWVVVx7Y3m830hkp24dfS4cVrH9
zErzNmXn5CqdMVAIuyizdE0aSFTLKlxHqEhkj8MPVV8n8Un/3M80rmqWcsG89UUbG6nogYcbrveW
t6T9AdWIG/cGBQl1bSmeIfdXUu0xwAe3zfnbgtCqGU8AVUuRfUu87hOsAlyvXS+R9dnldLLV/szy
SPggj+WwVGCEbIqg1lBxEonwY8GaJcyQTDWDfIti8NEeM3Ku5NkEGJHuf4aQBvkyGiKLW0BN0rSy
5Z3ZDJSJxpO3ZFaBpFYUqdWwG5v9es4nk+PBo5ceFrWlC5UVgeSwVC9wItws/FFLhBeD7UVxpycs
GgL3n1ZmHb/Szl+ymuOC5F8MAyawTlAjn+mgTPoT53M7RNdOnOd03aG8Gevpq7IAEfrj7Ma84lns
gejeqbg1BskatHEGhqAv/Tm9q3HdifpKefxZl31A5niW0T2vF1kOkaXHuqRM7a86Gjh76p3akQ0T
vI3opJHRZOcuGqnSjY6l9WlWT4KSf3QVEOR4s02D6RKgU7lRvL5q/HP5vSWeaCZVctnfK2JSXFPk
1qtXIdBjvlaZzkw0DM6nBC2nUGmEkXLeFvYnP2P5fV+6OI9MCihzvdYbAURoIv2B0HJ2cUdyKlgp
lPb4nvDdAIr8hndC9laO3T9SJfk2jhW7ER7tNgSTBzSbih9oedRsuM95FOz+mgZzQV9UpCi0K50N
jCS5pDNqRQRGvkveVmRGx38IM6/20SgMP5BeFnL7Mgpf6jCClxM3el9FNRf2RDw/10IXaMoMVl70
Xntl/5xNU8aWb2kvdqq7h+pwefSwPRuZLQE4GhOFZQTGdbF56D2JYgDU8X3GRC/t2tzuC90ctDHu
2cPJ1oTKlf5Gvh2hdW6WGTcIl0p06UQKtJ/pnuhNMvTIchqVGZR3UNCFHqYlXNnNLcX0TUFi1VML
CuePRprza6hwpRZwHHsRxwpFaXMugKNzfjQtpEgcqoEypauvLrlbNpLSQ58VdsAlPHtdTmJ131xQ
1PpAhD91ERDFElqX9s7rMc0EEgTBFmcXZrbshQj/ciiCQvlM+upzd9ZMf0pmLer9wk4sZVX/lFiw
5hUJwZgfqOrX5p49bkOyC4wiqkH53K9S6TL8bcX5l2GQg31f1DWoUG38FVRN3GpHzASfOJxCGr/v
VAaqG61sfVXz4l3JzG3r0sWhNkgQ1W3fuA2OXJAzkjjHybqp7K20FInQAxfYc9nsj6p0jVRewR0m
zInDHqfC1K/mx5H9EF/cGkIdiCfFg0Rr+4xFVQ2le/rbzkpum/8kk+EWkA3Or1OOvNBHDMbWQKBv
+8gwBgnI6YNQdmbOAM6KnDO+t8TWMQp5yv5c4rQIkl3bwsvg8vPsI9oPwbYiexVq8spopA5nv9xJ
dp9J52HEkgnN6IitAgmLT87uZhPUDDpBRZARJOpO32pzqJ5QSh2VNPOqsR1Z1QQj6JwTJt6baSEs
m4QChGpvEy4afpG/4DlfCGScBOeEfZUcBdvPRoh8lvgmiuYqXvhbcwK5evt8Fz67SNHSJGZAeqKR
07wq2vR0gcM9F5m5YtArPBvAIJMKPL+C8VzvI17zfKsEk5eMVg6CJHnFf57zsfJGJKeCC9CsamWE
5z4kzAb3sG3qM61uPbWSZL4h9Agha4ppUKJ4HjGLXnk/ANbbERjNk3T7A334R/YkfWmNhJSrn8oJ
90mf+j5apwTiXrSgTayDnmBjBW4tO7CkZQjc5KU9xaxifCZpYMYgHdXEL0rwYEr2WUNSz3m7vxyP
2hZ7JBs5dFBarEC0orLb2IxG5X3YdS9dKyi1Eor/r0oHe/46tB3JEpEDf/KbFG2ib7/ChjfBeKc0
nWHGA058+IwyqikXd2ujB0xLMldL4AnwU4mbbRJikZ/1OFoMcX5SjWBipBpULTG1ang4zXgBigeK
ttkjiblGdI/k+UFHCMQValyng2tdW6q5yYyUSc9rK24Sg4qgILHgle07JOGMdKSJHi2iKrGo7pAS
QcvMXIhH6EYf2najHhD9Idw8jORc0xvioebpZsyx3DWJ7FeI/2qxj6u2UIhBi/OslA36a+lCpabX
RtY7+ODoH2jN02by2Jh0xEoorTA3PzUJwoy8yMczBsyu3g6tnXzdxsy2TvOcDvWAeT5vwLHlDGyV
otz4cI2MOYQBHaSXJeAeNpG3yIRa/EuHKzeSoKBCQrgHNCJhKIY28d5uh7FlY1VM5ke7CiBpXcc1
UYsRyZTF5FrVcjd9Ke4L1c8XSlVv1GzJfRhf4UxQZXJa1yvI7tGcLaXK0fQwnkdX3LdY+ibJo/2H
UDn/sL2t8kU3K/jrGOTjRJyQzPtEsEU5/26vrX+KFkc0EU4rqQiT7lCv0E2Y+YKK2rMO6qLZ/CwA
d9TxJx6SqW1na7nk910dFJdP/hfYiPIseWc6/pFGUMSGpFSce70a4cGDVtUZs9ULIVErHsIPPFm2
j1hFAD1pojrQ32OjkTaKQSIO/8kMp8Gmtc/5IpkG24Dq5UyMLjBQhzSg84OepdPQ++5/atW0unU+
I+l1BDYQG9NqjSDWb0GlLYPYdEw0VTHvyqbZ8F6xm/J4M4uFaiM9M0enHRFVvYIDGC7LBcxhnvEI
KJ08Kwgdb7P/D4uAS55GC7bxgPQTN5YiHMXBawEIkIJ5eJENJgHPc+l7llm0GzatRWhoLgWZgv06
kUdqXN32gX4FPXtFobTLQZhkqJRasSvroxTPYmmKk9mtkDIY0ktuU04s86TsD6qgk3Zz7WwiEdcP
qZYry9vRmQvjANjfbKSHceK6kOtEY/2rsaHbQkPkhwjppf7ppNLVlsq4EfJ1gzRruEDTdxGToH5T
VWaH4vHb8z2uMZcqH5KQYUa2CVzUuTWAD1nn4cB3XTbeHaSZY/rnsHNxcGX5o2GccPc5YJZ6xByV
3pJxvjRvOszs1Ddv1eNBSf1F7z+IoqGQgvvkl/9BxHxFmtj3IDXBy8DFI4ENi3J883UY7jD1OQIs
uPkY+W+BKYLVJYLeLBwoEvgA/mWJz2cThPNslN5keXuftH+oGjG/PMf5s58BbkDJ7aAnvZ1SpvSv
x3uoYrh4E0j1SdJIu56hjGEXJ/azNrjYGPUYYT6e6btjjYoRss2mkyuBEFhPEILyrf3Qj8n/zkDF
fUhd4uE1i/IwBDGumBzsy2Gtt/KWbURdLJ222NntZi3ojl3sdnIJm04oBK7bNiarK6gBbaiRe+JE
1X47CajmK7eLUAqLTSPoQoJ7FZLR0gEfNs2x0zA9k0QwgM76ztPBsHT33WyhI3kfBrGa5h0HvEgG
o/ej1b/h2dilKybXLnc76QmzSXgiLL3MFdkfHz6QgpA3z70BsaE9XGH//MKTwsmzmklI8KDaWM4L
XDgYj0AdWrpRmp1EJav/9GsPc33OTmo6VXoFd8qh2JsZNWJdwoUxgeNnMDXPD6z6k0UV8qwVjHLV
NSg2HjNXpi+PCq2mwT4m0bVQDOAh0vpNSCKWt4TitaB/ZfK1YKGrLh6dLwXQMdx4oqiGt5uiSV5G
sm2IBUg9qgI5/y4S3hQ73KRxDKFGGcQkMuUkMsxicyk++EymTXtqc9QF3QDWTSnli27uWlZ+aIrZ
rn93tE8lAzl7EeFOFirUFspkezJ0/0bQoYNw7WhuiSl7J63RTZtwndp3jX+h8T0TbGftOu2pP3UG
X5m2aFiJIFkkjpGpfqVRpBPNL2N6Q60GBzy/gONLlWJFrFYtYzKsbm7ci1suFKte4HgeXhZwDfm+
ddytu2R3K6Kj4MJVl9btCMXm/srUmBiuUL+Q+3xv5eCzIjLzBsQdu59XFzFRkuUopamk6RDKRAuA
ysOyBDvN38pIqn1VjE1J2MUwnm+67ZpvURbLnpuUmlTg2YCgjaJRL1Vgleif/IcY61mQvCHxBgtO
BmnSGKiYmb2n8CxhMBBgb4KsU4J4D6CAlCaIOC4blWzdak7F7BuXzXp1lagcOoZg1oG60rahvXpQ
H/Y0SdbBOKUGsWyYv0sRsNUdTbwc6heubiLrklHuD0UiqW3s/T2DzQ5pRtaNTumGdjL6DEo86/iw
uE8puUYzkiTsBUvyBf4Z/4N8eU15tc5YX7d/gGXto2/2hfm0vzQKxgJNTEGgNSEAJTnvhYhakS5l
oFsJZ2amf3St6MYhtmbAVYDpGskiGs1Dbfivj+T89s91YCcpqgH6//DpZ+h+pc502OZhodCINgCZ
xqk+hs37bL1/kMGoTVSfEi4gywZ3VKqWUAm/LTrNhh6D9OHvQ9SBdFq7eJHrPKj1A+9bEprprD/U
+N1z4l6hOw6aLf/a9o9JMQ7IOeZo+7NadW21ngGcN4CnC/w/MrsvH2tjeq9bqTG5trf7R9UaS8Tc
5XOroOS3TxoP/EpDCYWfUhTYi8cWKrVY7+B0dRoDAShBaNGnsxwQpu72V9KbK2SzXgT2TmZTScNi
5BBqqMr5IXHwneNGRFC4UHWYNSgklXWdpGvPSL+Ty28wr+VOMx4RHgQfaQdshSg9tSfuYfn7mKWz
LqYqRsz2NiW9pxBZLC53irTtBGUayaKgeoRZXqKrg/DhY8QpcrfL+2glMUW22VOU5dHqY1QBbtuv
OnybX2AOa3Zea4wyJunhRm96m2ifu3z1cHBVpjwIYbpn653IDXphTh35gYSmmz9MrWol45kMMsW4
h1uJ9MLk0eIQFoVKDh8KRFd9uVZ+ugJmIpb68xv9Y2xp7UvIciIN0nFxs5fZM+3g7wrNzmYYzdXu
RNd0vpxerWPwFz74e4iJqLlJFmr0YPfPejUmYhTTIxLRxQps224B1lVY430Dc+jdlpxZHpTZVZ4Z
ziK9CClPti1KDyrWBnQZIDP/vjm/rh/wXI3IjWF+nHSV5LAEk/YgPpiRmNZX9lkBAXWhU3Qaw/xu
OOBx7ds3dOGz2Ov/wkHGwAi1ZpF/RVc30HaaRKzsqqzVfWAyA++1a0WfYV62qa4k9X6UIIkavcA/
/1d4sj+foudDfAZdN7PshCPTg71H8LqUEpYPwCvar210XSMC1WDWs91uzNqVDmJJCZ8MUf5TsjEP
ITI53ddTqYIsQgGryVRZXVF3VjzlOB7CAS+N+sEbAggCYicZ2JUZICQ//eFjPusgeEvHJroCfJZ4
MLCrdyQtqLeRnp+HVQNMe7ZIEpzYQQ5oElmfIxvM0opqE3Tw7PndPMsHKAPsV/dYsaIKRHa1dMqW
o2UhmHdBxM92iSuG/raG1QSsji/tzwtuzAbamKWJ3KYWGJDB1FcH1PzkdBpNEURmTZR7s6Hc3gku
OBCOb5qiRpr5ukUojV57YaCZYQk9iQoEp7Y8yNVLsz4uRMgB8E1u6TpcHqhj34dCo+HoZQhEVPV5
67mFEPiUEnHIVYOKx/Effy4dgQIv3uSO956j2xE67NOTYKyhyyd+WwqEiX/Y9KR3q66A6y3UyCo+
SFzh+PoeVcJ0sCInKgZHLn4hgVj2KNFYWdWu2MrFv2y5q67MkiUPHHSVyGde/IGPMWBxo8uDKduE
ExgbH3FbYl+IdxY6Z9s6PBYhIra73HTpyRYIKjiU8BaOkBYL3XhV9sfglS6OHiIV7RiBmSIinWJ1
CfBP/q9Z9h6RDXC3gEf4xprxDi075+urnHN7wBHEGnGxpiWWMlxcSXJGtTjBEt+vXx+L4E+LqWUe
GDR8LnNBgrF5H69OKPbezFs2y2zmXuS6OiRlm9/h1by9ze4iyWVoYTuKjL8/iW9GbOqMj6PwNV3c
BSXenreB8erp5jgYfKHouMMWzuSR/e3UA6yB6U4qMpGF9C1ceaigEGQp88exu947/IRo/8r7P4cm
i3M970UPXKGtjm6+wYZwmty1xBFoSQw8QYe1Tk8XsR7jx4n8v2RJsfbxpqGRHeuNdPKu7qBoy02V
mLs815ZTXjDVfW3pIJm1ZH4YG5tXTrFyr3QOt+Fdmz5TtXT6Iup2JoFdnQX+CekTYQpMg31f46RZ
9mwd8sD7dsFGdh4y6Zptq7D/sF8Qcz+SjuLSWGaRQ+pQ7MkKN9xHJPXLQ3JlBR7FQuW/RqCs5op3
4aVIij+m1C+IcUhdZUTuiHyvEOnMAO/16csc3u2meFUNgogOA3Bb1Yo9mhLizwoJgO08HVXl8enW
E2onQHmCZloRbUxYoDGkefKk2WvqrikM0Buz+iast7no/KB7zIrg8LsAQxPHw4sxtIBvZe8QY0rG
zfsV7Z5BNVdcGn/mA70fqLnT4zKa2mSirP7VfqgyyMHfCJzMU7bAUPy89sZoLb+eFs/2xnjLBV+h
hD4DBxgKHVCoRoTm+jY/c+6cp4HhEcdqpNS8grAZ81xBjmnGn36xkO3hV21dX7EwL/6NgPt2HiYQ
9PtPa4bpVhDzJNVeGbBeD2HgrPnpJEErAU7ayHsV4uWKgTn+M6o4KY3voqPMqCfxBnoQYwmsrrDp
imrdo18k5dZuOt59u9rDh1Yk/iouVJjTZUp24TY05elqzYAW8SaHLZiS+i+sBgWMFpEmR/2Sjos9
lOpPrd+wULeJAOuvw+oj8NJM0wD2r0N2PDd6wrmSe2YbQ8Tsqf7faeBceSO5vRBzflFBOf0ppGv3
4rsavAaCc0qAZl7SHmf82jvg+cwk+8J1cQfE63yDdyN1lyuVJyObLsinI33JpkyOFLrqIbPDV+9d
ogxMgN9BOaCmRfE88luVdYijNefy4BzBkJco6Iq6MYj5Q7VFRw7lz/wdI5xBO/nvSpxMD88L2kNq
qZplKB4skN3OxOSk1PQDswspbYD9JAlkPYgGQWnhu+4BCxRgvHJhajFhpBDFmgJLa/61MSJsBfBi
yfE5sKP9XkZoA+0CxuobA2XEAhskkV/0US99ru1FDMJw92xqBZOuTFWC9yuOYDGYWgF1nOKu3N/6
BwEo/TWQYRYeIUA5kUcr7q37AZBl+GRLtpxietNu6oXQHWmJCrXbooT69xBP1HHWrJE8FnNxk/h9
d08qtGkLn0KZaNhXixvU9XeDhFe79Jjy2YkvT0kkB/3BDFFaD1Yzx2IdTMjmetjMfyWAKcao4OaB
kAjj1A06e5W3e6BZ8HPiJ0Web/rWXA0nb/lQk4I+ATtgmxM0ilCF/f7kI4+f3nLK2X5Pl1mPQEEm
evP8hVn85Xv+lnL+34qCMUyZKkl9VzOn6GwAbR0zU3boqAz7Ly9GWDQ7LZ50y4FvME+u5ulB7KQH
jYem1n1qLMjc8GxLKsoJ8soKXZwcMBDVe0tEz1pNX8de6noem7RYUcg6YFnf4mtWuiFKiyHVHhYU
BqXeF4lp2KRChh019VHNHZn8dhebzBOG9F/7//griboa+Nma64Mf7GGRU2Qs8iULv1TbeBrNqoUg
kFxPWefIQwwxdjjpDsdYXUF6hoLE3WKI4uiIIMNXluOOFtD7S+9pnoR88fpDd4EHSqzuEvvUxTFT
8xIZPmT6J3hQFGz+oZnfNxfxlsBnfq/k17MPbSoO4hfedPJe/Vrt2ujzj8XjbHGf0b3c3GcDcMjc
lNjZhP/H6jrSnE8GizIh/4BATQlb2J1KD4ziy+c3ou8Q5nVOW9rI0A5NyTTv0jfPbC1Ojtf4M2oY
M4EILNGe42r5mPX+cjCGLWCCVBTLmtA8Z3oa3+w5mjZMFQYehnZxWrIHNWQ8ff3towifC+NAQRnu
syRcCjIbc6TPYy78XdY+De1+I6bKqLLvahSaKovt0Ng3j5flltSHNxsMn72X/nervpepbFiIVg/S
2PDU5UaQaYFrQMOsbJY5v1H1m62JJnJrEzIWZheEGeoTchkOpqIhBxb7d5/2+7kaES/Apl/kEABx
8E4bnHQGePkTyNdIhJy7ScboA7V35VFaGKUprHx7ZeTHFNJVtSuPpYCQZB8NXvjifpeqicWjnQNu
rx953NrL2/pPeyGtuzDYzAuUhMcvVhOk8bAYpMNdLKzGQ6f/0Y+sL6rz9a6KlULgTefuTulChj2e
bBz532vm1K4+8J76r8JFzJs/uX61Mx+ZQR2RKN0scEl2IQkN15inLzz2lMp40KuOZqJ+rJmh20N4
vW4Gdd8uSRoQMf1uNQDCbXyTgQj1vFvuAS3j5jmiIaHi8iejTdnveadGc8FWCIjITQoaP9uHynCR
cLEQge/vROogmxOxE1/hAmP6Ly0z/hRwsijK94BhJJRGGArwkqO+FD0ESxPAUzW6+LPA6AA+F7d9
HHB+FAeSjiPU4dVKzsenZHaoimSWYneAQfzuhnMIrA45mnI+iWWEPzym6IcJGI1eO7C+xJVLhoPg
dJFQ1olni0EgMyTuuFP7SEVjbyK4wlIxlv9jo4R8zwNaRhQueUSOCFANQ1NQEOvOsd+gFnoP2jCr
V0mFlpmo1MrU5Q6NR0zhItRFZFdmhTwZf4riAHlpmRU9KJfiUUPQNbtkEKCjsMlknV0PtgfhG5yv
Eja6Ku+vEbrE5pkplzk42WBaqJX2PLcmb+8zfEVkSu2j/LDkI1jhwIi9EFGX20h1JF1zIM9D6LTv
SEkX0rPaMtzUALjDexF/PJ74zMWW8uqA5pESD/MiblQvgQcSI2ntv91TuVXDyVc1t7SMtw4SyxvH
Q4AeSH2MgDFCJw0zsdNiBA0l8tyrqbtqlZt4DR5oEnYGE5BH53w1buJ13aYw3d9XYodefu1RXpVd
N0wuVFpEtyKQH6u118tbiDv/zDL9UtPJklqkJrrSky1QvWtdLdqaMcryNm91CrOA4dnivZ1lJPu/
l4rqcUXZ8TzXqB5Xbcmz8JnQ5PoiOv19Ek0+xpXdB7Ac1Sms4SrhPLUSQupdTr5saowdRxjds7GY
73F+zm3PNJOQhr0v75LBjpNHmFILvaO84t443I3Yq+t9Xylx3IJXz0wb8UrjFO52Yjt16cnTOACC
ubifjndXy0KPDfPUYWvZlTRq/uNtD+M/HSfS/pcoQuVghhfdTBFfP5BBT55D/RDLFIuUfJTJB8pQ
iWytL/PFk94dqBeGd0AnIkKfJTOV1FmL1dOXm4TkwVLy/RR8NzsT4IR/drzLRiMJ/SxJsY4Tdg8Z
HQjmgZcB1j+AR/3oCkyGvT7DxJGfYebMGiZMsfQTbk4676zS8bKnuHzNeAp8N3IS5KfiKcu02ut7
NIqtXrchD5yDAOjiZdYYh+LHq509ZJU6ANGMGdkBUIhLnwl8ePgGfLBs0jrFtqZodjkwm22H0G9/
doN+WSeBvt12tOV1FJPGq1sQQfLFUoZmG9dOUKPn5HEzS4rajg7JrNlh7C3WsPh6nFEloE2eW7iB
OMmBVkv81kRmk2YtB2e1Bf+BIM4syoEmSu633lY6+5LLCpbR246ghcNlfZaiP5qgk4iRm+ruk5Dj
2dY6hEd09ThJVwO4cs+Q1ozw0OZoVz3wrwjkc5HkOyaXGSQbguqbjpCSgYcvPM2KSiZb1zyTxder
wPN93G57ujqsVUip04ktfLpgtQPvYyZg2Dwkiw41G0uD8Tcs/E3WvZR3ZwRISopUEWFERHEmVdnp
/BTiExsHFZu1icr10uuYdMSVnLGdPSeXWFTmkyenDlnkyhWsMjrO0s54G18Jb8EPpUJKBfS83mqZ
SMrE7eL4NZ5VZzgTRxrZvrYlOMZ4MdnV9VUCroY3y1DhJQi0BwVMdWBQXuA190TW/+wuj1vyKBjM
NR+SgoAxr0nyR9cWgtTaUhoPEIFZ6DyT38UUKMRCycMqwPgSE95UNgRhU5fwxLtPfXxRpw5V14CW
T+e5eEOuMFMcqDZgmRYv0cNGhPsXunJCd62dBIkCPMSUtw+89aDkb2VEfh0Uzm6IMLOSjiGN8xi1
qjnlmmpGla2ryviMz+DH35aPXOjta+Evv76dM9AYDgO5vj4jm3PNR5jtoG74Y5TFmHoemya2MJGo
cMLT2EjCymRQAdMfoL1HpVGIYp9ShncPg0Inan27la3AwJYAsr5r7AwR40H/mawzMRBeec8SZFFc
H4zHVSYO6QfM+mieSL51niLGQT1FCVbV0BXsn03vRd73LBnpAIJYpjEthVOF7obYywDJe5KwaUPY
BoPU+t6H8cglRZfZkj0Bu0MfL34qOID7Xj7HEoHYyZLKGdXPoOqf8eJpntrZelWNNcho3cNcIi0t
UAT/Yt1dWChnPBr7BSUL/dLjND/jPca3ik2q1zelgtSvxSFfE/8+/wEk19OUMPKfqIIxjnBzl73/
EUgF+ODv7swShX3F2Uid8D/ym+j+NwyLa4LrshcQq5PFHppMvTs+ArEwPy895q2AxbTYPBMDMbqi
QQ+cSrSanL++T9ILrejpdjDx4u/zie4TRZLA4wTnBKn18vVOhUS8uu391fQRiSM8eMrj+ZApqtFI
h5O/dfSsjxcu0CpTaOAsVJdCpSF85g0XeAh1bmHHvqtdmo8JOOWFWZOOPErzmTkRpwJ94n18ldNi
IQcW5afxiOWXsUGsd+LjOpM7hjBVKrF6AwLbvhRhPxaCsUG7K/aPgPzjvmfVXdLBhQ6w4CYnhvt6
WDL2hvBWDs4MX408EnTTHnyZsfuWYyMiFjMbj4uCw89lRFzaQzibIfWhnRxo2xhvBoRjTXZRHcHs
HMxRaLaunC7YZW348jmz3UagRgaDxgUZNk5gu0y/Llk1kA1A+BgOGYCit8Lkc8Y4BF14pfugjcEB
YmnYEmbH9BrMTFsN9o8OT7uJ9FHC6NqkOXUaBjiVT8yw0wLtm2D0D+WzELB634A5G2J5wOVUWl7x
YKIlphzTzl2mGdYg8cZH/HgK3yN/W0RrpHNdDXKI1Y6/jNC3klHxzDwkW0pH9JwvgwM5pB+goVFF
q7SxyEUYXF1rITA/XDl/FqG13KsBHrh4//LzdjtyAiwtJtc7lO7IUhK22jyrDDxPDwwqI/NcrHRY
JmLN7b24zxKQh3kixT98e9tHNOdev/CxWyX2UtAav1mPXxa4NF0LP6GiH1ypz/zjc3rnohG3gT/x
dB7e5eTPZ3SgJGAvhJxt8h+kcLWaZ2ppV0GM9pQbT85yZ0XvaqVsKYZPvyrEK9tfLZ7ouhrv7R/M
RL1DV5en1YqseOK5ck1uSGBnvm1wskrUkpVrxYvEa+RY5kYcqMqTqpM1OK869hVzjGfmKCi5odCW
+iofVsJUG/LfYaoR91yamQK06KsTnbcfyK5Eemz7x/R7UrcrzS+o1Fkoqeji3OlkpGLz4ImwJqZA
DPeUOPVYo4eW472PbS5YifZSjfdJVmj8OpTGI0ee2/BdV0Uo6o5pDe6HIIQ2eBUA5jXUXF7HBwKb
EXzQQGDT6Znt1fD2FQeD5F/STaTaSltwZ0F2zt2ai3x/0s5i6tBG4e4Ea/EN1i/OgTX9DoxavpO6
9ABA5WAeXNO3f5OsBxJ1VYP3H8bQnA6UCoWqynDckho0IwuZdmX7nhi1RItL5eC0GKz5PzXoNAbz
4qJa4luO0RWWUNqYlQ6G8PWYUx70bLc7VY8ztquik+w4qFWPgd119lA9zLkFzCmibUWJUWninfOM
eBwQBcWwAB6sNRpzLkxLUMfFt3SmrL7vzts3HHrsdZhEFeGZamHup7zV9R8+KR00EQdbOemLVTyB
GOjlBkH/IYMovdxH9AinUeyjUMGNHW2qg7nKeuKANerPpRpCVZUqDiJZLdjHsKNVY0oJQ52sNNgm
CVpJ58QlPgAIVcxjrCCB4gFkWNitH5QGeGGE/H/k2UNJAx4aU4hl5t+ok4ok50jGwoVLCMf1lfgX
DY7OScD7oGfoI1+uJCXHT+zpdoMdI1YUyUc8Dkwta+sTbjewoEnULmKMX1ZivbOrKGf4WZLCi3wI
IAzIWxt5c1hm3vpkdZU7EgxbE4KQT0iDe7SaXOooTHWxMV7dkQRD7OdDguHZ6s8KDcLaUPXmhlHi
oNqvCmdbbMweF6FIo9/HZ+mpfF4qUT9BeXAjRW7fSKxdt3v0I+vOG6w/zjZJrxlYls4SuDL4WQBW
kw5ZDPkoDGNnDPMer1J59fa6msEjIspFJyAr3CQK4eWTfRvAiFPf6Sqd3byPUn5XMibr0C78M0V2
DBRfRCtyPag/3I9/GaSYmxbSgbGeAFe0Pg1l2MVjB98XQyYBz/GfSPxknqZpwmHDQS95xB6LCXy9
E4FG+ygpaA0ePZZr0Mhk6UiszI0OT4DT+0qZFNyb1Q2+vEVnMIp+a+H+wg0UJeuPmI3CKrjp+2i5
7DmuTEwujEKyu45LYaI0glL4S8lX7pees24yvgBCTMYUfXZbaHImztg6/wdOk48ye8WaEiCTGoC5
DLustXJ7Z5rWW2z6e/zpOdBZFuXXckRKIk1NAdWzbNEukwsP2w68UZDvio00S75xV8EqGCiT5zvC
MlNG6PGiIzn7kROfNANUKMh0/ycCDa4ZEOGG9mOgcufdihQmQf0qj9SGYb1MwC/O22d7poxoPlfz
OdxnnP4vxg58N5G9Yoix037kE007sGcq/YC20hvoZLRwThbq4d6vNaOFiinABJy22iS7VJVt7Z8l
gSe4gH3hyHNzTgBEG5ZcWXYaU1ZRLavRSPzJe9sCCsawo6M2/enIwOUVvlc27ZQzYgWpHmT25BdZ
7ZBUhIP3kO90yKwJUjASVS4Eg6TDlIuanF7YjAsOMb2MIfq/f3j7TjKA+vYl1P5AN5Aa9nyIDlDd
o6nwZUMJzDk2VAO6plZbHRoLSdbdf3eWp4g8f4zd2D4/ivz6mVJbjtvAEFfNdMXhSErXJ90IqWqJ
Kn+jUsFfmGwvD3PInQvAUn+4v5RGbVSbB/b06fZbnAEbs5YASId9INQURVWEB7aOnOJTWU12bYKM
fFNwEzCetueXxIlILiFAmX0mdyiC94bTU0znjFe1at3AAgzzs/NyX4jAPHNS2qQhKLdEP2AwuzeP
jYXeHSjNVjFP5X47cynjbVMs46JX4aoenU1qJ7BJ3j69qWy9LJcGla/Mn/bmDYSAIYXNpmHYxGPn
MvfhJ0llMj5rk/Krzr0hTBfHJGrjEcex764zGPBo27JHWG87vSv1WiFQVyJUPyE/GU7miILUTm4m
8U9dtOQkt8KSkTdnRbEiCwd8wgkrc/kR6cYqv5o6oQyzSo0Ft2dK0hjDyAl/V1QuWHMnEjxrj8gk
PDS1U4VU/BhCDFOfRGGGpHyhZFL/kzBewfWKKErtAnOXOvWzjZ+TqetVLYCoPShpDnFU89HVTD6m
J//Cf0o19o3Ul6bymGc5XYPDccQOhumpa3O4PLREQB7v8xXrQzOlHBkO9usrnuoZBhGf3zYMWafD
6z7rQ32MPBB3wnVhyd5D2yx3C1U1I0nx1NUngNvyszDS3Acv5YuX9u3P/x62sjKX0k/HVNaRI1w2
wmHW/nLdhuKFqeSDPb4P/zD22BrWPht+7rTNqghQG+dmomme7EQ+Xwh71Azl15w3WgsJcxFtJSyg
vhqarGGTLSdQpuq6SeexjJ1uBZWmbYPgTWRxJrGTxyORE/xfxHbU/rwAUly+Zjdd/N3Tk3VQF1q0
PD4R24HjTYaWw8HMO+7OZ4yg0bWVMylAjfu/cQsgk408pbc9vEFWQuL71ebGvT2sd5+gpap3wKdY
8U+BoNe3XCYoPqhX7FvYUlmyPJMNPHYl7tIwS24CsVsMmItwMaDww4fROmWLjkFMQYU0aAoQXPYZ
3pLDM0walrqUqfTq98A85fC2u4IdLwGqNu8JMVP6DzfCZVWLsTfpMOvzgh07+g5oJCaG/hNgFKMB
zbeb3GRDRYQuHnMcrT2JDRoRxUw87cRRPFunLxisg6NIrnP6PkyuqusY2DpiXaBg7RTve8z+GB38
XhiMbQbfqCtnZUEuaJ5Mj+/HeackwJx90GvZ31WLlq5NOjZ0SolY13u4MjfnoI9xPXCAqIzF/XBE
T4etCnIT1CS94F5e9XvzPKGg3eHxrCeIEzKpg+HVW9oEdF8CTS4hL7zGeYVMF5ioPnqse5EEzu++
lHdGEGkYODXVLwh78tjt6+3AOEg+AteUL40DEuTy8n0tfInU70VjXfVhVhd2JTZD7aRtfcCXcSeq
2z95V/zRIwqE6RHhdxs8341VV4XYGRuap8UKXBDj8ZIyHzI6GBemR/x6YOimGRTiI4spcUpw5GQU
TypiTDe3RBtW8CyCCnuS0PF0VCRzbe0R+/MAEOXgkt8m2DfAzBndPVQlbqAGB19m2poUhtBTcRWO
vpcBqk40KtTceooR33uEYMRlyRac9PZz1/lfEx4rXlHuA1JDTbhtVB7AeV6y7aZqI5Ocx39A50sH
bzQnLk7hVCEPV87hFDcc8OONPqxQUn7RbKryEIza2CIgclI3eeRu7APR22e125udDIF3SkkkbqhF
AGiZi5M6Ya21Si28gLYXli8OPlbXjyikiiRZw4rat5Bv9ESRHvXtWP1rUIfkJXmERiOsRnsSydwW
Vcwp8qmqkDyPUvdqnPs4vjvBzZh5XX053aYo0VjbuZ50llnexsSrBsaiRLIPztm4JhIWN6G0CXUT
vYTSIWpyHm9G9GGGdXKfJHxTdQL6AQRKrLiSAZHi1LMWAOEI41Dc1L7roVydKb4DMaLx80oIP4lm
k6xHivLE4hERErWfqjyqYYHEE52RpLChPmGksPC2Wf9pjIrX+wzfoSVanLPxUuCvZK1ff87Ny3Qb
4JYtbKxD30XTnSf7X3dKoSKNrAx9X50ugH4HGHa3Ltc6LawDPuJvb9onJT4SYJIQMSBXJE8l8gLH
TnpVA1p8W3tJcNp/Nwx33kqgffSsUQRhzKIoGHvd8FJqSdGve/+B+K/UIA8pdwS+dl5NJgvAYd0J
aa2+DMnRHLCVYcM7AshOMy73NjC6OQutMcEiLg90SiO57FCO70iGNmnfJQEJRmorQ5cU8w3wYJpf
04wTWMxX9UOhAzsXXtsP+bYlT2arsjnx4fQER82TaQYrOl1c2D4oFUmtYIwvOrX0lqB0rIpR9XfV
GXS62g1ylfY7TZbXaOrG0dYmgJd61AORAJrksLeHzPytrIJRiH5p/5yse2cp5mxLTTe6Kjih/Mmo
morkCgqs/L1sMliKif3eOr1oMHlory3inbVx3+dhet5nLFVwbje4eppSe/fkCnWUzASn9oL0a7Q8
BLVCQtljBlVbvXSASuPIDPFKEN3HOhRD5AMtPxrLlmGGAPja1PJoT1pNMTY+j/ROHrmazMWfHNuy
NF0Yulm28OSOsv1vd5T9mVOvv+RNImUVRQL/dbYe1bZHjYe4a1HCnPzzg2nwwI98vE33q2zd3CYz
KemsI9sBgdMsfecFTKpkD/M+GBvIIN6nhu7RHW/lOFevYHpSHcqj8tSGG3U0KaQC135Neshl/I/U
vZLJGOzRRk2JodDYdS7Bd/f340s7unmuL5jdFN7KapDkKyxjbCXjwUzTZ9aNfdrO/patC7jRSfhe
XvlptkVZkDgPwQRdKqLxx73gbxEUzmuEnlYEMww+nUefKbLvMGrjEMZiBagaWZQ1GzDMx54luaHN
7OpKNOwm6UcMus+/Ksb5wFTYZ69Z8Up3wkmtb2wIeHRSmiblZLWhMh/Ioh/9Fm9yApUmJN3uMUpX
zOiVhlOGSkfWNXKIcD6HOxVUnAH4b8RRXIxBEM6L6aLWaTEyaq8m6YWhs8it4ROc+B4n6UfjaOs0
BK6D5cmF6BU4Cj4uW6uaQ8QojxQX4Dy+k9qRQWe/WouUjuxBFnRrwzijF+VbVrXIctfgc2aNbocX
Dxk0g+wufh4Izi9wd4pTkWKeAs1lDQcREUqSJjIwGS8ipADsFEGjhLqb7ojfAz6j0pCdCfiHLP/I
COJEokSacMZnU2wyB9yOon8n5n0SCUOCq7NvDpWbD5x6BFH9smePL37VF5tHVXnmHFlpdq7MIBPG
bBvrWHWnfz1QGPp0K7qeJk+d3rGR8dtGME0Qk01rXe/OFwuNsLWoTLPvnlDzeInzSHL+7Y1OetJx
A5e9SXM8PqWRUSdZugM9PzdK6t75sb4yI+pPLIao+7AvlaHYeEXsQUn+ipNamQBO3F7GhS2kuRr0
0TSSdSGBOM+gbCECIbjOqOmAYJqpJ4sPwggzHZvwHGqALzNdxwdCY4pNsPIejke48X9ajJg9bBj/
aJFjo8qbntoL/jR+2/p9+wFL3lWs6jGbor5WCGbnMRa8MoUUSASLML9LWSGze9pW65BE+rSYJ9F7
JEbMPY/L+jRA/brNdtoyxLyiN4hySMLhxtbJXYsDV+N1Y5cTq1WH7y6D2a5fns75rlMIZjsPQtsI
g3ftl6WJ+cQLK+5BEcuzKsKK2yEsm3HaMVwKaNluHCnLU65UmYeNyg0AfgWSKz8Q5U+P+XDVWdPV
jRd+gU2jJr5o0PmkzPhNg+MBMjDMvLDV1/O4nAfY/qljHvwDyKf+vDsO/tB2Ld2XYc5xblMz2w+o
ho7JxcQIPx0mxwdQW4xYowOd/CtNT62he1oqIqIMNXJBBFAt+3KWdkO7v4rslPLlgxsZgoRGfVdP
5uCtQRz5NpFpiwdTS+hWG5O6CBteXI9fvSDX6mxRNDx1NUb1BUxwaNgivWhxBgKOp6Yn7F4wj+fn
Wj+VsoeexqpiEeMs3PMdtIRIXWSBy7heet14WQQEmZzEzzcM67seLcqNQJOX3Rb9dWjXrswUPxUR
8baDJdxrlZMEDau//WGixzKR9nQybc2kBgczeK3DDlYIkE/PXo4eSDGjKYEjiLpjNJ4T8NjplW1x
c7beHnBtDsCmXRk8ygHONZt+Jlj1etPybKXpUYxM8b+2tD0TDNOaNawzKrF4xusVcjsIVNSzIhJ+
/YH9ACWdk/6j+KUUNkUCpwcsbbPk9HJt3MYFFZ7tYbmk5vftrewUDlCo5LsIF2ylpu9cPKPXbOWV
XdgSUmLJY9wAsrnAVsvRuh93TpQgyfeQLcgQyxFJUCASU42D4aY6nO1UyN87QO9XkOrRd1xP0ctl
1vHf/B6Ad4hmUDe2RJX4lYJ+yNhq1xEhm5My+kt8NrK0qsoljDapEgVhv5TE25w1xsOeKhzepGTH
qHWNF1RTDEzuB92Eq0xzIUZLbHvhv+4UHUnlMvKU6iV26XZjCoByCD6jrCWLNgPuUBG29o3+X21F
Qj3akaOmk3jvvPTWhw0C3KMNV8ffuh+4q49pydMcwehUJ7HFzC8QYX9sBWLv6F3krCu7RwYASMMF
5SwGX5UNxzXuJQcVzp7PlwyagHr/JsuTr5j/0I9WcdGX0TqfNWyinoaMkAIDPt9V47bHUiek0HTc
o+jqEAJPWfyptGykaAnrCj5l7Py7Rh7Pv/56orSfMZOCGWPn/IjEepZjWd1Qv4ENqMVdbKlJ5Mkp
FE0Mj4MswapRot5atoRhcicq+l60xV2CVXymlF67Gx6IZLRcRSeTflyVZnII2+1f7wtXgGUkYDpz
Z/rm3IsB7khm8y+wj4Mxvgnkju/onyS57pthodWzSmC/edLz35r0PNKwrxrIvSaVGK04NGQkcTcr
Trbz9oDZi37Wfzz2HHxR+OjDTchdm1r1T9LHiqerStkbxwTP1tWSBBp1yxkEw8RXwwnIIiytb3+J
1XTDJDGJnY6cKfElGaHLhHXDi2k+OnkgBqjLGOmCWF4cgootgt9jdzbRdBjU9VUx36uNqEEgfwOU
J5Es16Zi5dx5leHRFvBL0b7tKRd12T17nD6TfJ8GgfseieOrqhrgOQq3Ipels+xm73PcS0IC9dnt
GzHnel39Q6K+y/VnYqqKjKwT8n4IHHpt6tLYcBILvYDzLgK/bsP1dI7z44QJDxbxcUgAAJngu8fT
5q6RBZyh/emkPvdvB/pIoTSQ8Sj8wRHm/Cuf/IPzSdsRc7kNVdxTEisdx2K0fKgv5kXfKQGvOXH6
rX6g0U7GHrZxXtb7g4RTdjaL6Ymm4n1m0I9nNxGyxSDFJzxLJ6lod2mLIrmv4Fhd64bkY5Mlm7DL
xOVU87vn8cLBqi90PdtVwKQRmm3rC1s/iI+XkTl7Gy+8NKmCdKdQyFOKTRsPryyUiRYAREFEJ104
I3tNmAPMrScAeiSbly2Mc2sZpxDCo63KevH8H9JcugHPo8b+5jW9yJUzDAQLyR4LBuyvRf1xQkyQ
/Yyfpl7enPPuF7cLdpta8m+4wBD/IKMDUxzrjiMh8SMA0CwRqq6uG9WCb2iPcSUubvA7S0Vltnlv
SU5+hSOQhwXbH8JjxNTrxYZk+3XoPRHWr3EgeINsSBhbG52kGVPqQ36/OXsLUURSdcjr6Xh7w8xQ
Xp4pKgk8huLgUMgQl1WUxHUr4ji227jFvCCy7VC2nmIytabs0qBkFW7yEDW9Pkux9z5Ih4tklpcw
pgI4yZnSHvGkEzZ8RrdSxMvUMzhfgmbShTBtIeb2y4I5ni4pFivQdsZC8nI585s8DJZIEN7z/ntI
OpwcwLGEU1yYs5srT1o5fSG6N9AfcLYF0vkQqhHSOmepunn+OLCQbu6eAfied42dKblcUTUoNsMa
Jg+v9/G4sLxAP4PFzTReMbdgRy1HS0Lue3VMBYyW2lTvjqSOwazZ12zQoxIWkOus1BFD12rTsgME
Nw6BGg2PrGyJaP/G3artxY98P2AwD8Wivkx0pow25sNqTKfKIek1zF+Jy5PrlyZASqVdok6Y3m+X
Oi6LQd43qGFP3CJH+FpO2W+YSpqPdcLuzAbvI+iEuym3vFYqpbV5h5XNA/DFjx93cvlgCmbMzlAE
bfB/JZ/sIIO2VbUmJdg+Du1vYSbtJGLul8AYMuy5iJeKk1Kd1IENWgX3G4OR1xpSupIAAjoZh/LD
obCjW1AKbHX3CyayilXzBjEc6fJj9A4khWcfgewM938PpnbirrwmvobSand1MNxpoJrogGLgWIde
DJ+h51eOWwZ/LcrbWQfSsgoodioS5jXfJS8ceYHANKjSMQITmnzdTinmiSv3TzLrpikUz9L/vpWf
Jo34S1VGTMdKxLuP8hOxeN+O+l+IDgIziQP0+moKHcEntxmXzfcX1WePjpTZMsorcxKmbFDn0aii
kToJhg6i5SADXXmVlvwfrShy0B9VDprrMnt04fuexUhXCoDagzAUeEUucjkmD0cUkiIxO472PhBt
5r2lTx8W7CJmP5ebUKELzIeedCaDVeTe09ri6VOMT8jFm4zJM2t1yrB2VcmcqH9UMNDrn7Q/pjng
0g95le/fve5G8wB1gkgVrI7iS19eOQZPq8gFr4vlpjxsDKhteBbp79blV3et8nuF1am2Rw/HMKMk
4DXNbQ8Q43LIH0578r/Y1B48Jj+NqTa+vM+bBgTCh8UjWBqP6D4y0n6V7N8stGIV+dt2vl/Yfiz1
/E4IwSeZ+uDaNArMpg8FvMr1/4snbIUeQCkLga8sfhSnuF9UO/QMKGkN+t7ImNpE6Cf/jJ520JZ0
A7lX17TtqbGTqqSmODKBcGh2j05HvHS5OJhQ2b3krnSrh5tUS4tGXy70sOZjSyms0oY/VWsHXFHC
z9mHhTJhWxIr1tB9nHgaCqXMmlzdKZohywzL/QzklJzKYFPajuslolkuFj6r0mXzYCukkFqminxu
GkPHArjKEQZx8JsKc9aFjinguDlX2nG2YPJE9nSlJoNd/74LrlkgqTxDDXC2UHPlCKXZzlNA3PK8
/w+paFa/qD+hmXk7eQD9H41HPhiEqQdi4m3H1rJnhqHzIW8eGytJAveabuBip+E6kmgWqq4gznjB
pfAnT/+94TtkeQEoz65/YSsUyFMKg+CnULfOQXnE1c1inJpEVX7I50uk+HQj9HRNkFXM9HXMNE9P
lqG9ib8pV15QHuHvVSpBcFjYmmtYuMrq4L6RZnKZqDsBRe+4caMfss6jYoUynEJbD6oug/XuSpBq
OwxdsDB/Cajk8qbu5AkUh43GEffPb8+GRbXmRPnS1vgoV5FIfjSMzGNG4hIkhgl/OMloQWKzEYVv
rMp8+w/0bnHWI2VxH837Tc0CWVWxwvArnpT5QvfvmyKD6w65WrS4n0EJxqCq8fIHJUt1fhjchX4J
oXxaREtsdD6Wv/GLOyePmHwJ72g5M/S/aD0PS6Uh+GeKBYqBpFcg+tjBCkn+LDKv7k49DBRY3rhn
dCdyNVIgOxOfnBylqtxnGlUkDhj1fPEC9DQtu81O93xoNajvtxrYsBCrtcH3Q/53EUV76vDB7oWn
ZtQFmL0GZghVLxeZimTmnnMrhYeMy0VtCBLk+PQyZBZWq3TNoebiI4plNyuEGiBi1m3XZ+1jlkmE
ITI2NJ5J8zUbazb0z3+QlRoW3eEZky4lqQ8AZ3gEnRa4L9GqghMs5gpKSi09kipVAvHCnH+vGEbd
qvf+soOjDVUTLIQ2IJKvGjVlZQPwwD2JO0xaNyNPK3EsJ5ZufJfM3UNUSXE4sxUMs4Sj97pYOff6
8aBxElPI3JYU57Bt29zZKmLIX1zQft6m28OX4b3fVWLJwUgF4JocJg5OKmfDKttcIMgrGmm770cN
O0HRG/Nz6uB03NKyiXAyytbRLi/OU+krJsVXG1SP9VF7n8pdGFnW6Zg+jF1LNfiChD5BAplKAJNC
ebBihS3aIboswhobu4ZR0qmVNvUu8ybSPT5zTjGFKilphNzVZo0O5CUqIEBep1cWkhxe+GXXZrmq
UXbTQ8BUZV4ron1xaXD+k+GFo3d3dFY/L1UAnGTmpNFaYWjlJwbUv3iKdEWXDLjeaxKsbwvb8NQw
p4M4n09/kLELh7wXgYB0Y9o5obxdRQQHIV2RSza3JA1R7rS4aK+0tjcfSPuf3dqXYq9LsSLTucTB
qmsLnBPyM2YQI40F5cTdZua0e9Z5ORE1X2l0maj5Pp0ML7GcLHo5qSaD3Jaw6DEHK1tm2eLkaXEK
iH3CjUe8wl2uNeNiAHn1kfSeiWm1jYVzTLPJ2E7U9ODa7yd7lGGVTSZL4CsvZJfXRdAetZbQA6oz
/iqcpz7146MRXtkQgR55A81lZjBUBg8h4cXmkqxFDyAOpmIbGQz3SXMswPd77k0W702Js9gAPbVf
br+FC6cyGvHDDn4UCteCuPRM3dZotUNlFFxGh/5Ai/2bcaCie1fcy4gAwuaZvQhAMoyqwnLQSvCw
v30ZtJwetPzmhhWj2pLFnkrkmJV3Vu/Gj74sl2GGlp/5Cdw8gmsuEDNhx6NdAVJDqUC4RcaPznUy
MLaZceZXyZc6QLxqBsB+TnJl7nSdoDdR4bQdc5zyZtQ2H9WcNZDrsYgxPItk6BobigZPlKSu1sVH
tjyoH+U/Cg74S7CJvWWUWBImTgtEzD91axMHUaci0SoRp20BuYjuQr/8UYN+so36iiuTW7f/P7I2
ELsk4vN0IdkgrId/SmGZBwXKpaYm9Agb5JHQzACE3uvKQ7xxFoofqN2EfWI1lLdEPG2idFAoCAPp
wtTGbSHOQoD1fdQZDdTw8jweEcMxflwmEvFDieGDPMG4Od6VnSHl+TmUeSncdoi3E1PrrOElj1VR
31L1cTgnrxLaIvAOoTSTrnKDD1W8KuTIved79uH0FPfDeIxGGFNCPikLY3CS2pBatX7LKm84mTcc
W5bXABTl3YFNCGXUDJ4/RQI+TByr/d0j6aqtuJpufGsR7y+cKLnQV7p+8TJSkUtw8z2pqhmEPrh7
yO0RUgNce4LqZDr8ZSSo7YF2Uq16URmVMUHWhSFV1643bxO/uoWab6NKuWC4btT8MomAONtGVTz3
474Fcv+30f16KwG764HRlgllypE7AZo1oqPNgVcwqHcmluHe2ZW1tQ0kXqFE99t+Y0YzxHCf44HT
/DXn81zKVsCwcbCnr+uJcIDhznH+4+xpW9lK6S8iijJtLq5378rC8kB+dzBapc5iR+YfSgO/FkAW
Hc+vvq70rKLb6vET1BVvhCZn3xAIlxdUSg1b19R+ZP0eDDlt/cB+pQdM0HFJ0Xln/isHEwnvodrR
yV6bTLfhPEYnbhlbMnWvFFarquSe8Uux1X65Nnj23g2Hi9nR7hL5bm3BW+e9s+0vXKRWXqqC2P38
umuCTgmRcelgbDUGZWwRx0wNExjshjnaGehhXjAROcqG9jOe/pPaM8oXR5rsINlzlB6ETzFnYrDA
2q736LTPHOnaNbh25nikqbACfaoMRE4iUx3qVZjakv/aZ0yrCr5ZV9LFdWWmvGT2fkUm5BORYsTF
fewdlgO4aBVPMkzdzQHWRpV+pLxYMu9w38OuRiMN0rPFV7GRDckR6CGRbKtnvNO9mr1UjqRVcXRk
8nVwTxc1tZkCO523UhxI702Ym9PiYKkXUwUvcPUXUuG0us0fbePsiuDf+hDw7BFnnL88rSjYsVNW
cL4XKLgr3QXqdE5ail/S6hOpdLiFbWAkwKVQSPJ4NKxVcu1TwNDoZ5bkwOAI/QSO5Hrsb6BUhakD
9Q1VH5lY/Vu31JVByj0+tOOEqtuP+YdL6Fu48Qq6BXhtXr/tDvdqJHy84bpqKnaeHALh/ocwJ7HP
xbodgkAPb+6CF/hv29U+kMb+0u5NzSMXA19PDqsGNZBW2aI3/Q/Jr6XE89RFGPXruBj9jR/Oq/cP
RaSyini8puSdyQ3Y9+p/acQP68aw/pUcJoZrnBmCnvF8YE41eoTikUyiJfvD9iHsesK1nYfZN0lc
1//pZ+nC3cfmB2V3uvgfML3TYG/B9CZOtouy9RlySmRqEtW1kWddFYtMUHCPw+wg6dYzeDsCe7VS
glUzhgrIvGyNOjOJHFylLB2FbrsOOreEkjDJeZnCjMB7fBWu/UIAUQ8z2u1B3cmykAJH6bMmNTAp
3CtH8yRfobFxavGAFs00xMJwUPkve+4J+gt7cWwmU1kQxdMab+3SwQ9ClAhlM8WZyP5aHX6ERguS
UGD4+cKabWdErYqgsWE/YXu7ZGPPFqXJmvBFyDr4ldI7IBuPWtNPOcQbKQtEiqdVDZkkOK/ew5CE
X54rAXtJ4bgeFatcZvx/5obFYpJH0ng+OCCC4d4cPSbIrZGxwo/0Za5NLMk4Dt6j5TeubP1lV62W
t2fpUQlJS067nAEtXRylPdvcvvzq6IAaQNHnmBZFCKfa9Nckruum4UW24JHvLjH5I7prAP7s7ppy
tpAMELORmyg3wfnYSoftB4gMCLNSkWyEnozb/+fpbEfvI+dVyGVg3pQJ7hntLUnr7xjzWRJGjPcO
gap+iFQunND3Q0Em/K2RrwIaw+KDyuyeGTJGzhrEjZo+agRDN1gVZTav/cG/HEflkD/l/k2gOKgx
fARUF4Uci2E49SicsylMEIzffu56mxv2rdg1Cjy+B2L9byFkVSbBdXhLricLC1QkBEgD5IH+m5lm
HujsMEhzB6HjQedzvWXUp3biftSB7mrQfRFkxP9EsfqbgKkxNnZ4F9XVlt764KoHnFkBVT9TfzOj
O+LnkmcweNDj7YGeIKT+jwOe9iNhTd15vlMcVnDTOvQ11ExzEs0MmcILOOTI8Y/xOevhKp1u5+h8
jr1GXtyD0qGmV/iXt3qYvEvHnxapQd96yImR6IEoHijruv5/cewF9kf6Pw7jIiFUD19Oc5HLDtDh
aCUeRaQuktvBW4T2VdHhpElwgPkkrr5xzezjC389NMMcDSKhgxl7E8XXQzaBGex40JvFVakK7Tj9
FzY3a9Bz7v57Y+9jwFE5Tpwt4uFSeJTr7iieJw+UwWPqHY0jDF5FOMVUs9QCJgf4HnWlnjTfbRnY
dSvVerxYgqLHtusdJXveGYn4HR/LMogFQCQV5Ew30cT3YhJqdYhpbs2Pv30nEsuO+nzPb0o6OkXg
B7i6FTdm9dII98USFRcVV/YIUetS8S9cz8VNck/ugsK7+prNof1QgpgWz0W2YRZ+u8q4wlE7Apa4
u4lAHG5sdvx1Bi0r0/kzQQ4eH1ACfntzdE4DMSRw5Wg+xfr3mthBT1l9T6VErrQQuVX5Rq1MQPgY
Dvmdcex5iFBncwT1NGuf9HCSxokLgFcwjCPws3Xn2W2+4BRBlV/TZQU1UpztTHRehnvWsCVTGiUt
oK+LJx+nUvPV89QB0NTSvP8mg6qggsJNzdfX3B3U8SviG2FXaVnIAuT6iCBYIWhjuf7bgWaiAqQn
giHPrNz6ge8BcQUPxEDG1Tf1+4e6pF+PatKE1O0w8BPNk9AtF7jsJiLntxL7CJ3z/Uj+nV3amb12
carVo0chChEcewQ3+0f71pCY+Q+x9g8MuMXGIzLWDlplLKM/n2Zsvn74FzhYSodTvHGVIVIYqGCN
VNLCfNW4lgzfp2mKqbD3Cp4c+rvZNOmZqTdcw6vooUUdih/ztkQ+2eAN69dt5dpTfefqMNqvliJl
+kp7R8I2rfXRzXhuuqguDr59u9y4CF70tHzCG3MFg7qdu1wUVOB5hv3ZhlxWOm6bIhyTHBcR3Pya
ocMngK47F7rz8DS0YT8zqO6L+HdmWgJ7htvMzl/kgL3HIGuBUGXdvH3m3eDDjjcy2FqmNhnU3Lsb
g8JWtYy0/0CDGdnSeJuiVgepRgLUQSNgPuOP4aPUocjUL/PpP8YHbq+rdcmd0GECs7K5WsRVmsES
M3cxy5NTeNYqBqtoEgGqxSxkV+i8ny3Wzn0nbamRyhp4WNg+7e+m8AuvKmYA6KSjV3B6DnIkzi99
mE4CTQEw+rQhr9vu/BTgzCtgun1d8M1KnM15BP3F6dA2PTHyhKwrAPayB7wNEU0u3d1zRgjkMcud
TEAw2tBSAMrfXzH+9XUIr0DQgKePImcAlc8tQqVWraFptPLDFcj9oWTqqW+F4yBRNQ/GJEECEdE/
QgPXq1AXrn0xNtVqAkNWeVTlT828f319QpsggCHq9wIFKjhOCq/PM+x85JehnLnwVkI+NudOr0mH
AnhU7pLvwF+KjShp0pFw5z+7grQa9qfjZj4PeX5YdfBK7N7CyXYqtMJBdGkVP9qPiRmgGoWSjxAG
c1jTeanpyFPRrd5ftTJ9gJ4k0QYPrNHfbwN0q45LluHZK4ntGfPAuBWuBwej8hTv1ecL0AqEaJb5
v5qDP8SxZxwbGnJDEtIvsoC6CAKt+oxnLPDetwwWD6Nyu3UWoBV4Np6P0WUJ7P7Fp619IbtLmo9B
AEA09AhyOZjW+DO+g4xyIIV9Q4la/4hyS45DrxCAn+VsinBqrCLB5D3ClC9mgf0yKZYOFRP+H/Sp
LcGUjIrwImKWEstlr0X8oIEm+wvC9gbsNLD16mYaYfVBhg3DLspqo2BlKw6UK2MBf8NZKqScJTgd
deQI+YqnCFLpNu041WlEdztMHWfg9BroK151pZLIa6Gkpe6T3CmA1FAK0SJSka6R9maIzskpGfu2
J0mH2P1bMPCFJXYFNF2xKd0mvxOqqmufjMgdtl1yO0/v6yYT03GwLUybOKSb3Q035VjM1zV90fq5
ef4G38iMHBw97bDuoTP2xpb9EH3KiNKtjkp7obv7mC9tIQ00kdOWGyHXbBg9BkmwDG5fp6lGYzFc
/WsS02FG3Pl405Hqr/msslyuQQX9cdnEnPFvShEq1KLs44iKBhXEBsY5/BAgXZ+BujAkOM4zeJ88
azJZTCn+9Lh9YeQnVgqNNJ/MA+HnSMzgijfj0q1+l4ENynN0k6xmUjmtlRyEkSQjBzvMGxFTvBTi
I+AqRsP1f+wjrDXTidoAYsRBHMeZgRKtwDKRXg4Bpf0CDga04Kc6CXBrQHFkWsGgWy7fae+kkdO6
CPs94t96x0TMgKsM3f9i3p9scLD0+NScbpT26z0zpomy2zCf2WtT5yJk/rjCaFjFsd4AdrxNfvr8
osTAAR12pl+/QtwfBIzgg+sS3JhKvzS8xKnvVbflBPfRrbOxPWs0n6rJDszArY7D6SvC9tJhy5Hy
IYXm9nj9EfeCpgOppLR3vgTeMpaHO415jGgw30rW8PozAEqzPTfzlzRGEdhWpiwjyTIYUbLcXsPu
aNxxxsf8tfe6TBywaWAy8gXxGQvSR43nSkjLAUYNHiXQHMoxUc2/Z4+a9BiNgG2Al8DZIJAgiNlM
y+4ITZukUXW32myJ3G3uqRLAKAsaMNQt25/1nmGMvqPPpqRmyq9ZHAGE+Gzdy7aZnSFJERrFB0si
Buv682Mo1QJ8YCfQMCXTVouuDKHfjtP5o9A1cAx4hQmG5vL/pwluFwP2D+JQc/HAYrkOOnTVidUY
gfNPAJ07xaEzbAAXYevBMf+NLPKpjZ2asFyym3FVXnutgnboAZiGtwGX/4MoAgr8C8xPonZzDUlc
Mrjie8rqhk+Vly0bVZA/uGrixcaLIBBFIND7Ca9Hry0TliVM9Va0DrtR2hwvXERdiR0ze2xGSqXM
8U9H+fOUvLDcEI7xXYbLg7aXmUcp1hBHkrftlHhb1ZhOmnbXOw2S2S8BxoCSpilfF5NdkruR6DUY
7r67z3UMhzymigSWrmCFa8EQ1nVGHY1dCPUhDtuWWsTNakhJup1ciubqHvzlsD3Ttp/dx+jDwJAP
Kd6Sr0IqvODhnb4Og1KWPBR5sckDnXV/H+7J8yw2KhTBdrSTapIUU/W3rNfp+d80pLlzXF14pVxn
NCC9GpDcEZ4ecxEtxzxuSEKbz/v3jSvSR143d4aR9/PhI0oiTi6PZaIvvtmFzJF6uHbmAjb1u6si
S26y4qkoeWQTOLpXt7Pnzb2jlw93VQvvT6qxwIOqahc6N3M7Izle0uBoC7AvmTtVMsbiatoGWpeD
DwxSOUKoHXYnPMszhOfi23yVr674b5Euvg2VARz+5p78NeKgrHWo1LbvV7xxjH9FYaWGj5urA1Zu
0D4wJbUtIeTJDd6hNIv8paArBDeTwhmfh3/QdhXAcwaapkcfkx8opfwygKf0pXeNgVnsB2Rik3Zf
NkF0spPVcbC+jD2NMEqscdk6WEBpWsvPMsgKlfXo+xawOd9m0gITpWNpgfA0UaYUWo89A1ZUUsI0
4009YXzYgXhDXOBBC4zCkpw5xNxNtWcRqtK50F6W8WpsoF2hM1p6oFKhD3ptdA4RjODVpY/Hq/sW
PzELGcibxNpIBV5UHZkVWOxCwlajaVQKGufxHScioGQeKjbG6ooyzxzmZP8J7iBu/ofy3l2hOMRW
RikZcR4zOGKRVknruYwRZ0U5zBgRNEAP+e3KZDSldfdkufiZulcFG0JZBMs8rW7eiW0m5JIuzQIv
iZJNVIsUQyiExCh5nqLvG7DhiV4uYypM3GSEYNvkaijAQaQ3cHCzNtVPNZYjfgGcE4B/TEV0PT52
nRGadugurPO0i1CWH2v9nZAW3+XgpoFVP6KaIq1Z6i0WuLZs7JbCzEBifMyJX+xKy5xY5JJDvzTh
ZzRszkB7AHb/kVmRQkYYWGqPt6guKyTZ+ajRiciCDXxiNSuKTHdqLBHS8gXsXcPst7IaucBbxpXh
XMQnLcPP2J9Li3wNhM1OwtT0Hiabxx6P0yjYf9lPxADyA/Pj6Pg3/fMQw8UOWF8k4ms7malUiF+S
3PaaaO+zXVJ4GWxvB/gyW8zRTkxYrByrvyqvkyaB1kCRq17V2h5A44NELyG4OVQK5e0sKrgUm1Kz
JaYyQmIrd/MH2KyWh6IW0D2OFKrhPT3WGkBSVc8nRDwvJmbJs9e6LndToJE7TWLgU9Fu1ZGOTZHf
2tCeWCV2KMCnHLrunibTgEbU1BpAJhhD+V5tXx/1/TgzIyAOoNZKkE1MTH+ThySwSbo/35WII3G8
H4lsPngrFNNGqcIr8XyZmt0/8fmQ8KEdqykBzspxMjSyWh3KfcCl3vWtScGDoBb6pyGlMy9bpKat
ChyQS8EQmWgU0ryCL3kkXnk9OD5BTpojaGtYmHH42FA+mrzIOEuMPtq+e6HLy1Ex54B8YQCef2Gp
5uLGjtXIegHz0RF3Jl4E6ns1KFdd7DGKMyIMUhxiFsjiJ3lWZVyEwcmbUfzc7GxCyzknFiRBWvaZ
pVXXM89P2Y7tSDPAvsXtSmmlfWLWXESIwb/1x0zUme+RX8/3hahX2yxBFNt8ugqfc/VhcpjGpBWi
RCxeds0EY7Prd+o8Mx+IDrkp2Jf7hjy0+BqIK1+z7Z1XwcP5tFVlBDDrvL/wBcFFSPP4sRy3bw88
o8rmmPhUi9n/ypu3Nz1yMwvvFTFaYdKx2H6CKCLL3C3uEGPyVoNcAoJtW0gK58b7APc0h+hnzf/D
/XLxM0efs4U0czwVnUOXOPVgTA0WFdTdus6k0JXG2fTLU2oX+j3ECFaLlkEmlXYmSVDkbue0//vU
H+S5dM3avmYv2wSMzuZ0exRaB3olJ5S9GJh1VjzFcWU0dcX4o+9s2okIzvgp+gwTgbVzYD6cBlSO
MTGwOHvetCJwS9HZVZG8Cu3hobdgQSa9vLwkFm4OToP1Ax0ABeRUR74mHR9A+hE9RRSFB8WDlN0w
Zhh/7xqGhyMb9NU/7aan4jW2QHSZzrnAno38lbklywSNDpOOgEFpOBPlB5XTAsa7UPQBcMLDhGtX
r7MnNc7FmVePuJu7Adcnhg7Fye1F9kARXEwsjPynRBTSk6365B2FodsWn1n5b6xVNacuPHfMQPmA
esbDp0N52kCkqC6nTivX+swFbN+ZzD9H4eRZHVbW0/PgP6nq2BMjD8gtrreK0pHrXZBjMl8Ejr37
6Tzq8fBSBORzau1fs8lNHBph3Rf8MNIFnydjimGzoyNkwyLdXuHnqCKMFVTC7oMhNcSrL8t8NinI
lAytGR82PUXBMfqsfubmzqYKIR2YcxIsxzEQfvCmkQDKTC/94TGsr/nq8yNmoAIG/8ihBEk82orO
d8vPFP99d2eWqHrRAZAMk7FIxMjt0p6FRXCxpxvB5ghqU/DSM0W8tGmnnAuV8Bl3nL1FsazIeSqY
1FijqDdosaTiMmpg7uZVlo/unkkSfOOXCh2sDm1nc6xWB/lw+FuXDE9ivw0rEpKdT8cB0UMQch/B
NdbhmSMoeFI/uXjcbfu6Ilxd+MGMuqVsvNVdJWnFwek8v4ywGCUNHlzAYO8sRt9We1HH8XRec/lk
BjU0aJwoufgCE5xz0yCYV4dTV0xW88ydBGdP7eiiuD+SaqsAcD6uLBLaIQ/+9eqEkzs9265XvLXJ
/e5sSDBiaEB1ZS5wnjg0Pemyibb04MbD2Z5Rlw6w1kVoA0tJysSTzntlem7vTpQCw35EaHbbWFae
KOT+LI3s8nxFtbbJHtyUiyH4fukxVa6Eqr1dlPEm2LdNu0H6Ac7Zclqy2G2JpbeKX31ijjsDnQ8H
FXJEefb+gGEOejmLMaV91f00DgT3ExBH/v7MIrJs9bT5bw/hWXimHMxD33iCRMNHNgKoVaRL1C/Z
CgnLCRd/GglRvtwfNaMvzrAY0z5ws49a/Z1sI43iQy+YdMi9QBkWQCuplIepQ+RFgdkmppVVvtnW
jq3PGGmApFL1ZIkiqbIm2vDXHMZXCiV/jPzlxo6UKCBG95ZCKnGuLA/w2vyO3HKQCZMv8XcGnXKC
hlgDf0Tp/7Ftb/p0sGT7jTb+swSSqFhEfvlSVnTF9R8GnZqx8Ub9tXHb0FR9PjFJzEtfCCxMe0gF
7NpuQOmdULJXN799Etwq9UWBivsI6XOgaeEo5zfLjidii5IGWKIQnyz1BjcG9huZpr6B/gCpIoSH
xg2ZRIj0LHN2X068VzojH++slYqz6/fIho8GQp8rseIinU/e3VjMiDBJZ9Ln/tj/XfTWON6oywNg
VAXFnrNY3qyQirnwZQ2hCeHjaUpWn8Rdsz0/v5TTR0NWmEnx/Z4wqv+j2sEzklav4Ac3O4OFxbFs
I8CxX9ssvd+k1eh+cyfOoourTtIQBFG3RaGICs7RTSkr02RM74OhefUM00jxP10ejvRfDBF5i4An
zl6AUUfI8N6TcbU0K9TduQ6epizoOt/s4S9cjpOJjZlFia5A3LeFpTmpjb0Jqj2b0whSVi8wR1hs
4BqeZsgLjgrd5L7Ztl9bOa5iaCwrPXPWzy6Kq/oE8GID2ivsY5Kjpolw3AKVKQIstrKJacJVY5xH
urqQG3v+4Zzdjr/OWMHL0wj+RE/Tb0H8Cmbaug7wWXwBrbVP1nJxBoFlu6qkGdN6R6RpdSMbZf6Z
R8yuxG1FoXiRDbRV0mbF1iqAkP1E9q9Q5j6rV1T/5Dv9uj36UYp3rdqxFoXB7ZUhmUyot8od1bJ9
JSEXT1Onu3hTb09IwFXDlkPsShGZD7EXwoaCAIxrC0LKUS/DmRprE6e7rOCw9HpO3RJ3RdW4/4um
xKkBfmw0g757/CKeVlr38Gt84DpEnuzvPPUUfvzeHb/FjuEjwrblt2OviiSQZ7M8qDG68wFpYbR3
MutERhclDF/vxF8aGb07HtZfi+xSISoRX4skweqaOZSf+Fqf+TRZ8x7f+X24NjjpMj9VoO1fYezn
I76B3hOwAbW4zonLlj/JcnNjZe/z2yRWpQ1nJrHfS7rb0ZVb1+t5eElqe4DfOKBQWiYA3W/kQVjk
tZ1374cXbwANl80FJFMr+hk9z+D7IvPA2wYsNnUzoSOpQYo/O4ea6opP/wFgmlfpZy4ASh6hX8yo
ioRMYnxwz7SaKohl163OSxkgN6vnFYn5yIHaMLF6Cy+ErzYGELSgSBUDOb1q+7z5l6W8FnonHfmv
w9UeD1Nf5lK87x07OJF78yfnNIJYiaJX4y1o/aE/PTau84PsUf10AXulebrH5Ua6p/fwugsK5Wt9
Rt+/BefwgRA3+wE47OIgsJg7ut+ki/GfuhaZ3SrtjtSWwR5W8gD/ZppbsgjypoSR6pJRz0STDlJU
STrWhRD/r7CQhS7fN5ly3t9il6LPq/oNl8TA2pvBw/ioplwI30ES71VUQUkhMeLn1OMa3P0aWdYL
H/IHMEEiEHHWqGFWdsqdA8OKrIX7G/DEb9V028ZGKVv1P7jgNmS0FXb9uiWYGyD46WEzACTOIeCy
lSJkXGELADu60Gdc8l+KU9criYgYYkQK0SkcUp9AFZDsTvBgti5meVTV2TM99vY2LMcT3zjxBS0t
Vt1dFIVhNALUgT/oWiUSJ3eUjakD8TnAXbfWbyM7fK9z+69+GvfYnTvqgIt/QCdQAYDqQrREFaQ7
4amo/kHEnMnAF6YQZ0tROTKJtHeUXNULxUn4ONtJefX1NHCleFVXAHlzgR1o2L5TgpoAPJ/KDw7I
7L5cdNbEhjw5GZkBrnTlvc9NF7TZdobmAQrja5s0wP5LhB8vScNwt1ULj0n6SzftABz7r7Yaj1WJ
nqyHWdA5L8DxzrOgc4FC8iOT2fLVx+0hYVtJ0a+qndZ+SMwE66gsZ48GDtarF9Kpa1heEImF3vWE
Dmsm5A01uCSsrvazHYJZTDylrVEGbLRwMW3UW4vyBsUO3HWRzl1lMgbgbN/CDt19JY1GLZInON98
XyQ0H7elUKZiKI44HBuFFBwLD7uuMRfXctFFM4I/DnD9F1ZqGnESeRTQHcVIu7+o9crDIxj9A4Iu
vdVlCNK28vwCqKTSgEWPhbjV9hUQukxoIpKzuu6x0vxCtfYSZ5NQzg3cKrBSTQPnkKepOG3nlG21
THcTBoRAlE3eCqbXOg/U4ujwW1l1Vxh+wx1TcxUQ44eQRKYIVpauzyq6r2sniHVG1V4K0a1ddoko
qdTAqbGWLFEm2AH48i0F5ZY1Ivd+xccn5cmz6d2DveWHAB6behLa6knbpwJBXcWh6ASLhpRnhW1I
Q8iSxHmiKaJhq6WlmRusaAe51rPcCNqYS1nXvuZIxD1GGNFgsDRGFCgADKgzfMQ5owz62MQJno+b
h19eO8rMAyD8NCpI4TMQ08VuePMTbjlNC0ftQ2SH5Aog8Woj7WRCF/GFniCh4VYO86asDOHD0hhH
FhaSQ2JqAY1TVDcfpr1U9EyXYgG/1tERHUGIfVODnCvc0zum6DSIotn96aI8RLaQY4RaHo6dbGqZ
WhUFj5BoP1001zqGkV+i24GTI8oAER5lLo8zklxWOFKT1fY9yzJoztE18kW3fJaTPcGHP1iVS5CT
B5IeGzzswhdJ6OFd/tBhpBpeS+dhiIAzAWoMJfwoVTBHnZFUfP4dHOqz8RgXRw41yj/+DM7j+XTy
bmd4oQzfqOgerEsi6A+fF9Z7AnR6ebhjcuEVpgd6c63XiQ9iyvq3EjhqNpgHq+W6MnlxObkLX/j1
c4qciBFSa93du9nq5dWsTSLAmWIqDtE8YcqKgFcpDJJ34q/sL4Un1SlUFVrIvgQ+Miw6Ev64OkH/
cQsiz+Xocv+Q7GW3yHqdl1da9t+Q8OE36ot5bOkHPItSOmu5OOEBDK9oATxS56+ZD1+6YsaZl5aX
UA0kCs7Q6DOBkj6/+vlCnjGiIWFiWMJ0Q5tP9Udy+cePdRXi5ioIxkWhzwOJu6R16V1+I64VplDh
qleEYwHBuNK/6TLfpZG/6s2tzg+8VqUaS8cdDnLaaMTCTelLVMxr/nmue8Wp460ac3cpkkZVE4yQ
CpIoTT0cSipfu1oSSzUut3K10vzTUU/+QovuLRBbLmdyLDQ/F+rPiQgFMXYpHz/LNUgOEQm7jTAH
V6ntaBWcp1MdzRmz1D0ng9HIT8ZeVd22VPLv1EBqemkfYq7oF9zPmzD0viq6nibQ34aRKOHAAoZT
0ZFnD0xUxFClq9pzPoN+qdWWhjk2ygW0GMZhWBnz4BTKIZU040iZRF0I8e2lDu9LP+zuUcZFBW5k
m3+oM8KOL7Vr+XUzbIG4LusoT/g7e8LneofAy9v49yMLZCzBWQBbt5zXwqP+RizNCBzs4Qjc6mXz
docbxtX09SWJaoSsoOfhLVI1o6zVmI6IqTRjAdQWALTyuD1Ovp004ZqXSMtFjaFA+W7r1msBj3ZS
5Rs5e+Ut20t9ieIQC7cwk2nY8SXwY17P4r3Y8y7ECEZN2vVea9yx3nm+uDmfBe5J1RcF1pWJr3Jm
AGExPmOgCkiya1sj7nQnivgXUfYG5NHSs0fEPtghTng3/LrbRg718UlCJrVg2oUEuG63w9+paLjQ
vaIyIqAa9/BEeHoYVG6FbxU9PhIIMOanBStpVjwuZRBHJ8BSS1PPcF1VKvalZWE/eO8YPvMF509w
/CI2iH+31M9TV5LwhXUwSIF3LzPqvH5JYsW3XNbsTRciDk2rlAJkkcaARXK4QoxGWGjwOqwmU6DC
4zY+czHejPVim6m7YvZ63kmG6bKJkAK8vb1mQ4zDXFqfDhhAMMx2bYKVCGkCoLnFTFJ82igYnNee
OWr/1SyJVzpWJoDm74ZpajYrRzMsl2MAVe9eYjR9DdiNMYVQ8Nmo75mx5jVj1H4hV6dxW95EO6xj
dxHwbykkc1R8ivcxDazt4+YqVDZW8fRFdvcRebp1KYLONXEhOqYZWupayuZsT4TuO2iZqiLDS5rA
n/9VvSEVJzh9XhfT3xhft/Uas8pAo+yZkskYGYMq4U2EFVegaVDWn4vB5p6D1tJBs3s4D1Acomqr
5d0ToEKiwPidjJXLQ7q7ZgLzga3hXeqoEHfNIyLvdNk7ladm3MB/Wjw493dLCTDsvorZs3FLlSLt
zO0/ofpeRxtxNz6yHKl/xlUfUQwP3W+eMt9cLCl2maksXaC9wqonNfrJ8zdqh6tE8VAu6kin48x+
Rrylk0KdQHqu3dJYMOkdVBYFak5IxlQeXdFaqVLyCj355D8HddGZQmaGI0gKI8U/bUWs+CaTIOB1
UynBezvAoOcUWZwhBhWzjo5l1Vkie5s5qwmQPdi7dVGmJPLjQNVahZ5NZbp+G+UgAqET0+jBaRFQ
zP2H649myl7a38DKgI4dpbgs4hbZC9x7NGZUK/uvQj6EvdJdY7ymzNku3VRseGnpoxbCbFkO8Z0b
MUqN9CQGA6ID33frmGVCXNc4QVAu+72umC2k2QDQ6c9cde0JnuJkOCahOLT6y5oHK8/qyxxGWibN
DvSTSHclyXCP3AA3vvIgmnXC2iAie1wRh3EOefsC3RHPlMFtzYdhuV4COBcn0i6wGQ9HUFWnf8er
RbBnDV1GVnlUxRb/IUDWAvb2sXtqCXr5rYxumSvzEtYLiWFaTgPh+3YmQLBGXlxq+QGLkcbn/qyc
BLiEsfZs4vANaXmoAeg7iWr3ASSDSibizLCXw27Lt2jieWmmMHLnIIvmCY8gSamzGFGxiLP1OKBb
nA3o37A4OTi+PGzP6TLuVaVNsILXpZvmPrJnOgSXzc53kBKU5NmKctSvQaEX2TdcfU99N193wkwt
oaHe8EPMHnvDe4ycYYU/+vsp3woRFdbmaGgsvNz/Fcj/SqKLEZ5waS28ZrQrXx5ZD2nBxhJn179U
ar4oSNZw5eLagNZpCl/zvz2elc+Bv3Q0YGDlk8s4SqCrtLgfQ9zYUU5er/tM/gGNubkG/ub7f4cE
7X5BVtSeQsLekmkRz/kcN45cdA/XADON1F8MYftrSyzDnTyyYEcgksv2zMynWJ8hvsjy/LAjabuY
xn8wttEBxECmc+DoZ0ssbaJWXt0nJlYgBATgtBCqyAn0Nno1YTr9A5P7vtkoOMmtk9VnM4FCosv/
tfNwjpfAr8uW58/9tU6A8BW4qk82Jjz4CTuH2/rcCZPqziUVP52Tgx/LLi7/Zk6nZurm8q6JgeMe
TBJBUIsUstoy4Lp/Rfw7FNCOu0YapEsF0YVjhO91UuL7wlS3ehOJXR+81pcF4Yi2V6BloK0lU3rN
K4429oK6IAieL7RhUq/Sj9zE+lRzvexIHZp9RTjYjF16ArK8SL7VmfMPH/TOE5upHyRad0dKyV5z
35hPSt2cpCfgqoeHmbKfUtVoZyRPX3zrFHY3VuQtcEmMwxp6nrgQ3SAaXdUwcV9AtNLGgh0T35RD
3zVRpRy5Nnk81hxUhH3rwVvpOH95OjdBbvFgNbW1OxCZE+096bxrS9UBv/SBkZr/b4PKZXp4BAhc
xei/C4iWIa9qvbQn2JQLCPsFTaE6Uv/rgXIsBoPrXMB3BuPiHJFvTv6nLVWCDILhCM7LNG2EuiT8
MeKF2ArRFlPZdLFbT66hF9lqkP3Dp1+JmuOTeG5+y/yYBE4FGud/s3TviH9jS+kMyuf8/Qe5kL2X
pvG5elV2t0P9/ddZty5gTSM/brOpPK88OkLYaO9x1oKZZ5DMsbD8m/mRETfmFe9Q5Fhc/363v2Or
9wsIvahS7nTbc/xXcgdszJtczxGKMQToa0Zg3yE29IKSLlXroXeSKgkqMDY3DnaDQ8OZfrY2DWlh
Tcakikk97LvdA5mIT7jtW2MYJd/eZyb4/RD/Qspf7wfav1ebl5UJwPI293U31P8KgjWZfTp90Szm
Up5xvsfnQpw/kyf0M2+IS9JT7jXih1ZOiv+UiXanZdHeKoIq3w0hEs5YprSnT0+Zrua/FI43mmtl
0a9mm8xOos4yhwtpd9ehYN+hqbYmyPDIbNmKGJ8fglaK7O1/YsQ+clo++GJaptFM9gRKN2wSpqja
QHaBxIukUXcGpRnXKU047ucL6g5TvQcZ00UAFNbiU0vXp4k24X9pn00oqwEW7TFEv3A6iZ9UQeRT
7QdZwCDb81oZpMjM64MTmqJakiHZlPFbT52SxxR/6fR2X83a08KXEd+bbZkZuJ6YLQmH+P/cgj1j
+ZMrQRFs2lIeFQ6IWVlM1epTcBkbo/tO7Oodr4DlwKWe7Ycq8sS1e/MXuCpim524WoIBlJ1QFllx
htG1+y4p4msPAbb3YQ3hZtxyYcq1ld8XtIE7UjlaC5pEN1GaDUi2vzOPLC9jsNGeqW7GjWA/gkYD
E+tCSPLlcuMEC/okmEBHKVOnOJ/skHKl6uSXii1X0oe1zK9Zg4FdsTpq1DI/unV2+lL6D9ONESY1
YF55H0mFMjCrnSgs/+0q43nIqb8+Gy2y4NeZsm5cUJzGlRufQdBcmnQ4e30los9KHL8SSlFHl8f4
wP0WBwQrWnD+j6cnhf6eSv1EDYSovRFv7+0/BH58TL96oVtc4envABUxdnmNwXv4zP2HOxWoR6ZL
lbZ0RxwCJ0uX/zKdGEOgRUFQbvcwJv72IZ0U6kpF/fj1vxZLaFUgyh6B8NLlGA8VDLL/0lLcTz5c
UNwT8Fj195b3sXjEiq5k33jxJJIXq3PTTcyWrWiaJ+Pa1sq/kJMh0qXQnXIm9mL4hPwMznQkjltO
cIZ7da9cMLH6CCEho5I1l3PHBs5ZLu9m0BsP6tbIe9iIP5RzndvMDKXTuIWsMglRAx+Mnr7rEymY
cB6V7P9XsEbL+Wo7WF9DoMke2n0sRY/f9Zu1iA2hCxbfAeAJUPjJehJYUPR2l1X8AOyHo5Losm0M
Env8agYYX6ExkqW0Cv3i6E4pmNMtov5TC0VHxJ3VdpHhn65wn+rCLP3RDHFpszLFLM8uiVmr9oal
vm/J6qo2hhQImJ9kn3Ft1bwDPYG2F+wjRW9KvRZzHL9kynQGm2x7dZv9RD3g8gV+CyC2s5GnVhVj
s3KMJ6MEClyBNc/S6vVDScJC5ihY/S8UiiAg06felYQWZs3MY8tnFQZaSQrWF6YM1kehx5J+X8WH
UDX0I28YwuzNZ4mMBdVLFs9BDvGBfMM7Sf8rlESIVVMZ8pM0Ntp1Rfih+y2+6goN6PMZy6/9q1NZ
iCGusMFi3TQcUbKIUIx1Er2yqwjm7fMRZfympJ2IDttsgmP+wnZBHYfrGBCl3Dh+Wi+HZJ7ZgZxm
P9rnONfF0rlLfVN6rBXDdcWbEnMKRm4ZiziJuAeMwQMwK3Dym8NATwQlJBt+2g8h434SoNHI7VDA
1mLqzira/zamYtraPrFlFnFodXXhu+1fcD//131+ZyygWuErDvrVcgXzhbj+SZbQjLt1D7jSlJOd
Ca9EnSoeE+4o6hnXg1EOKEuRmJZRrkgHzlQdg4gFa0urpVzqQkRMXCIG1yX3ZrFrLTxcHH1Mqi1b
0jKFRGIpCWsG4wq14S4IV5nwBRj3zO7P005m+q31RLKGHtlM4EETOcoYYUyY0WMbM3IYYh3Lo2L0
LdAvO/tMVEgOI7g+I53ZF+HcndUeVcxU9HX3thzYV112s8nfjT5IgKXlW28hJi4ECvocOaymDggG
VY85pd3ixUJenuQWDSpLyPwSQxPZpYFWfJJEkA2mYXmVS/PGyNWXTHJ693G9OnrO83oIMLzKgxp5
fLBAXYOPEPmDzIPdKas0Q7j6ORX1nKQaiUwEwogaXkqXf/8IU8Fn0oE/JKUlAzUMwJHLHaiKRpJ4
M2aCGLPft8AJX9r0Dm3u0N1TeYqDjQwYkVRWHIHPM6IKhmhGfTAjXJdl6UVEp6f/9o07NKXOtK5z
57iGSIRGO2RWNr3Jdevx+2551svEv85LG9skLd3R+ZbTzxQiv3+KdmVC2GWOOvbbGwFe+vIrVbSi
W+6oqQ2cCmGIKJ6XdYqQlLpT4k5K9s7k9Vn08V0gBGluA/nHFJinQq68TpD+EoNqVTpd+Ri92wQB
RA8UoLNinkDIIx20g/47H8uoV4xD+G0g29bSPB90A5340IQe1/N832hxcdCEG3lzNhvssYOB1Wdh
kum5zDJdOHGCdwcnGET7NRiVV/FOmTQhWCLCaG7o3EtObseeYC4jf9ZL2feDXyaAc9erH4fASU28
v2KnIxZ+HSQoNSYUQntO1JEtqWx/XHnTx6JOtF7VpQC9cMnz1jlFWnqixO19/uoBSKB0vwrRE5zw
YGkcXe1gU8ZDil9LlLcTtVoVJmVEBqDtGiAwaFvP6iS8GlXRutHfnjCYWfDIJiGgSOzzjOi9aj9Y
u/20pvyYHG92U1baL1PPUnf3bT0WgmP1DKOeM0nMLGzhacj1wlkLOux04tqJysLUkDkz0Fy5bcLR
Yf9WgfAPDsE1QzrPvmSph/mGPfpvhljiL63QR6zjrMAggFh2L/fJkPoiw19+dJ2w6Wu7fyQWV5/j
r0SRVQxR/p0OFp6GjlaCW+UOLgVCjAq7v4d6s0BwQtBRF7aaOMd5u0SFYoDIUlZZvnX3yirn0HNS
blgttHXKo7Go6fpm3S2iQmmpJBYLO+lPOdGV3FoMN1iB/AURD4+guZY1saI/tou8zLccCKdfc/xd
iqdgB3rxPQL6zKjVVccF0lZlzJoeQAgJ3wtdcM0pZrU/1cVlV/6o9ViyaeMO+PjvVSPweGe/cesq
8hvT2/Obj5s1eosnWkHIBS4YHPSKsPkJb71oBEYFSm6jbf8uQUTuqP8xUC9FoSi2cGQ4MAnu6Q9P
GzUbXD8ey/nelhEfAWha5DnGTpzB5q1rF3azdvhtX5x1sWyqybH0kfJ4guYHiOdEZbp9N5bmZ14u
PHBd+p8Z/b1y3DRJobns6QoobQnWLtC+Mq/KbG8brr+ZWvcebfCHTRdNAO67EUFqbKVVsxYLId2b
RjfPrxXXXHTk2M7gaPgdzL6faIl1n3GckxnIveTVIAuucJJ4TLH7BxjXzlDSVeIjwHiVPD5BuCuJ
Hn/agXS+W75cSRGSR2KINQ/l5Auc0DwHHQx/xbvl2G1lyiP5EdMlCeCfPfXtlb2LUs9Md5Q/i7wg
xfnSA8gkpfuIenlmWFABjdcrUySil0Ksdh5di2A0DFEffM6aitrk4ghkU1EofV7dc1xaJXlrj2V3
CqlvLJG8MDr8TpJaiBQ4qQ+Owb0x3euchOM4Fx1dLBhHSSZQT3uGXLezYk6pZuxELHDVoV83CxfW
YT30s0geOkm5GHe+9rBx8F87Px1zs2DDndVUjDsuM0OToOsYFmPiSuQh4q2mt7R6tRq+dGY+kWe7
d8I5opAqKlCZmZzXxzWMP9t6mQS5Xql4jJQ6ro9eHFX9QD+P9FyoUqvgyWvc0TPZKbyJkv1j8bH0
VEGzQ94SdvI0TNpz+X4pKuklzXffDyUEjifoTRtfzA9MxTZViSnhdn4YvgNm2TTFil0KvuIna8e9
p1S2mDmv3z2dMjyTwvi9FI+wgms7RRbZLacsNpU5aDHX37AusptIOohIS/c+uAsTnYFh3SCeX3Ue
rcE2209s44AChDmTcvoFwvOZ+sMhGGTIUGy9jNTe3X52kDTCU6UvrwZs7D/7/BkWDtuFykc1DTH+
TPMek6+gTsbwQIA8tuw32xLmQmNN/lb4te0o8f8hlaO5f3HWG7wS94clJJBJJhpQ9U45cssZFZ6H
5CnTaBFvvIPt0vEHePiUmhTEzfeUm+K61YtXoGkmQyVH6z3SGw5dQNX56UcGp6KJJUH+lP5PdhEu
WTDhck1Jfqsi6Snt+Duqw+jxOFMOlBXRCZkpjho823mLLkcOOQgj+P8wq2+klVAiKDXhD73A13JX
oUNPrdp3rr8mDpXYB15DKRANi/+YjIqVViYi7APN69WGizdoxETpROrwRsFTPSunXyWMdrmVI1GU
RdXmQOfTeflTXyWH7HEqLHCCD+LzjAYeAcEdPegMlaSYIqzGFH08UDhXObe1kjWud/L5LsWshkT7
dpZA5IYRjfaP4Zipj9vrbpn1vK9UswInOSXyzzO8iAldmNq723cwQil+OmMhJq6EZ1cnKf8BxDcj
XiaROTXwiKVIsCfQnKBZJautCshH7R14j9ZXR4f2q19zucwFqdnnOZ5xT0IwBnRVb1G8056UPx9h
KUl3hAL5HL1/s+RALWhyJAFw4gnVxrn365qOkG2B1Hk+nVPG9euz8PVYAoQG/tvE+ojoXq9/BFpB
n1bjkZ62KDMDPshJrBi9Xpw4NOndTbGP+0XIsxc7twpchuLH8XVkd1GnkxhTrAw5CTE97AZrnxGf
Ah3lCA64VenClqka5+fHnBV/wahEU6riVl3kqhyIijnC932/aaHtUyJw8swVM5+FrWsg38/uzNhc
pLkewt+hZ5FSTtLjKHWr6eAcO7EykgUToMWIUvKZAGBMUvyDgO/GHZkcluG2AQ7a/7xnun6MpveS
XnmQPMm0p4y9mVUAa3fahizW1viFlqERx/BqW2mryg94lypoK/x2O0ST7+sBOQl6jEq8Zqw1F7UF
gpLbWBbuqUWuwpb3gy2VMlbE+xOUe1gIqYcFeAfry5Ord9qEVXewtU042fbybw4sGWxr5b/TrJc8
/yAg0TD4hdeOyJIK8wHZhSZ7riaV554GnSTyzEanoJwVpP2jNVpbPHHQD/s286usTWFYEEZy7pwX
9zD5ytX6itnzwIQr8n76j9sO3rVcoC9P0BCaX4YWgwaUCBrAW57mMDrrYVvhQYEAGd5ZgQ5FFr7P
i8ge0/YslJDNx3/ub9wfzOpngFAoTwxFg7bvzty2L8V/9nl7EgnQQOOwks0JXBj7UhRYyySQCFEO
8DLKejH5B2vg8bzJXaSOlDeKwU1qiSOKhBqJ+/h5e0GCnKaAsMdsCtUvudwfw2t87t/r1gxKRqrd
7QMlcGJeetrZd4xNi/ykAt6biVWNIXxnqQyyP5vvLLDvW0ydjBs1WribBcGR5KNT8TyMTxEiJhsp
gXeC/a5lGlosl4+8F82ftuamwtgi4aNGwdRAL84KDhjVPmxxxHixLve6vAERjVxEXRL1eyUuxpzK
ExMpaJhuAJfGGJuYQ4JkCOf1BQHmKOKzLqUnA3zlh8Mnkj2MKYhermTadB4+n1RAoubkEF/RdZr6
S17WGithDGqU3cR1EQ0fdNGbGAhXnSV3Vt/FqgUsgPEuUlGcecdOi/pb4kAMnn9ZCfCpS04itWXT
617TVKdbRzZg6IsNAlpMPLZ3duVCHa2oHHT/WE8RVW4I0Q4k1isQcYy6o4qCMW1oCimu7tUou7As
CU7NNINeAVOBxUx+fVRmA/jN22eXa0bOjClQfX61SAMyaEPQWm/7Fcl1iNndpybouNeOH5ipHHhY
FvoswgDtIFIsmoIDyQnxBudXiUrCJjA/fAE+6mJcNQoQHnHfbGDqu+hZBBE8RgDtm+z2XMEVWSV/
s6nyjPF6fSeoY93yuQXMMWqjtXFQMsy+23DLLLHexemVgrG6/ZvzDKGNL0ZeDHpQQoUAMyf0LrW7
CpE7aWUyEcSZuzyRrVzAvKQvlvP5vPOOgXFjKu76Q+JIGHQk4zJqoqxZYkrAGuhbJ545awPXFWWB
hka8vThSOdK0c8T+P6XIyyZMW+Hxp05+IY4ztBK9+3cRi6J47Cuj7iffk5dfoPl7hHERyqyS3xKh
+arPqcZzQZgHACkd69eHAqdpOCVEI9b4DqWYswAO0iVjXEos0vtn+sVIAMzmABj2a7NLV+a+UUjq
/dZEqs4EWCfqZV3WmlL78zFNfJuLLcZ7gRxUEux93gxp8mz1tam6O2EpOw4EqfPs/uTpeuIvrNuN
dDYKfaw1L1RFdf/uQwtriMe17HfE0lAn5FldtAbP2NS+3bzxB3tXdX+trWnlG21y42OyoD3OjprX
EeBfcrQW1mQKERNyDeDMMMpvqFZy8M/nn69rrkrvBfuEl2meJ5GGMGc912GEOFL+yWLHkty2aFdn
SOZY6LGRzX2AMpG6v9N6KsQQhpaXIyBvrImUWBylzty8n4ICO8ye1DBUJ2hPRmi9xpr8217PXUjU
ZrlRQI4RUyJJCexj6NkSfYfPADXVQ99OnRKE1T6eUftY1FUF03EclCaweFbk95Lj2OcfY1V06hd8
uuooEfPZ8K+HBEH8qYFLfQeEq862/GOsoBhaoiYHC6kPvvO2vJ4soZTI7Em50cs+3Q94PslM5sG4
oYdMgxjQHzpwh4AHDb4SBY2aIwGC2jk+VMLlxLCtCrOJJ900vMR00JuceEapPdZTrN1t1gJ9zTT+
p6CAuy84fDVTVbU6wllzbygcSFY8aDBAo7Eb7OSS5ck1cuOFTCw2CO6yPdVoqaHnC4od9hXGgNXW
DFMk3FPjyKH6AZEGUvQmELRTYe8BgygWzwiFWSU3Hh+IcxQTOBdtc2tiNT6VaHxLI0rnGGkCeMoV
mDTyjQ55oT9j4JOhgYh6uKoviuSCcQHCGSTRHx9/hljYTt931RpxNpqn8lGGtJtnZD/PCZUsLnXl
PhtgwukgMzWKP8cSgBC9kDAAly+3TI1PFGEZPB9cO8TSGapMNHPouJ0aHOFkIVvrlYF0Qaf5TAUG
gqvnvItern26DonJ2uBV7NNbGLTk72vEvSbuINqtPdmKuGWatJYj6lQF8FsaweXAcaXtCPGuz41y
eznnoazlupLERB8mOm1dEuhG1KwCjpwDQD0AZn89NysHgH4gdSt9O9kya+f7CIXO8EBeo5JZchBd
fk8ykleizJQMxmk84wuAgqcGj6JO4wAW9RSfp0sSo3ae0Gn1WINLnSBDNir/KKHEA6PN72lMu0Wd
FBzddQLYHEG6SM4geFLdRew6QeaHuGeb3H+1Obvtya67Oo2hHl2t8XZa3hoWJfNlG4ifvuZCYT5f
dBcQWvvDdu1u+dvI8uH5PdbfKNguX7+xsJK/r5iLAKkRU4XYjYbCnHiIqVR8FkkGqn0/+2/rbOje
c6oHnIUe4hqDNjRcagefie4p1yeRKnrt4uQ6Myi9CCDYOe2JuF7s3CMNDR+wsZJwnx+YY5VocsS0
Fk+rz5CqAXNDoeunUkSYcdKOyDwOpUKTDe4x6O70sww47krFIzgI1jXSx+uPqFOIHiBvE+/EWkFD
cydwHI8SDVqba6sVuB3WCRL+yzrvBvatAa/FN0hN1yoib1VEci5zSoBnV94IwdDkIj15nWyHFXZX
omHbaGK229pnySx/SdaZVUklUyWnTgkgk0vh79cbuhUDwXXCe2PrWu6tLNQvBgihteDoJ78udx1E
x4V7rBL43KacJv9Si2tXRNEpd2XaHih/5GkrmgbQXUTh6xlR31ru8ZShuEvVH0ioqXrKfX1XTABe
ZVENyvdg4c8YEZYKWXoko1NvrdFch3lJhye1nPEE1iqGPzZcLqA0ei8QfYaAybVeZJ8tLYNT96OJ
OdSuTdBrvn7H6p19h6QX11ecyYc9ADEttmCbspJafrldxC2uP17Lr5yaSy4AqksLlogKpXUlYVeo
9AnmIXrq5Wn6qXtaSCwc9ze6mrfH6MaKFzy49aIkRYeoz5UFSitwPqbZ7yTYvU/V3xU0AUsQ0KgI
Fsgq+k8PR2MoLmrywaubdH9QWsf0yU9mBQHe83xh4sU5W45XQKuEtM0iTnn+lJ2MlteqVkqdiWti
uvHylcq/J+PhizvoCrS3ClrBs+yDBkzc3hh3ViOt6eGE/1GzmwNggpitcPHE4yaT5iPMEyjbTzui
TraPcfJEhroncuB375VREkpuHjqPydz9xem4S7y4aeASvOBe7RL+L6xQzMJyh7t7qG4WspgPAgi3
PhUOojxmjvlCU/TIJMP+lzrutAMeeYvkCcUKxYDB3MR1/EEn13i0CnhjFpg0dETrgD4stu2F5hRA
vx+RdrPbIJhhxHJqe+I4mHC1kPYsfatf/2zTVNJJflBCdxUtmHcbCiZRj+WIVh6w69hoQtZ0josn
WqrcT8gPCEUm1zHXpgT05pGNSW2u+2+f365ZOXg1bf2389xuXqBIc+nUXJNFqW0Ea8FZakIhmqjQ
lc1DSoYKBoHrttnXb8G8K7qFa1H2wRDP3XZ4fIGYX3EST4pTZVlM2tfSS95jlqVy0SIt+0CuTKiN
bqaOyOoTtLiL2XnbkE2OSp/+Hy2y++IdJnLBwfsZDIMmo/ULQblF1jDaqzxyFlPiJl51gncqXPul
khfhOeRECGX5BgHFp7bNWyq9CQTJsmf55vSOOjwnzzYyQScBDQMmVwdHTvDmJ6ldKL3Ftx1Q8d49
PgEsSOPvWGoDy/jz7kBBkLluLeUPfJj7PPIJynKyY61aOvGQ4XLBf5Ps85dlivMlf4uHE+LcsmHf
tU0t3KlAtMffX5puPT8+W4MsxWCzipQQcQx9fBy9dBtAFyl09Ca9XBduSgD9hyEibPt344bro2+l
Wmdw59cmjKt3aoI4sKoBo3Zn/oQrV7P6I42xSdyC6UbPmDfV497TVABD/AmLkyXf3yoPlB047cOG
DQEZfOQd/aTewXYl0BV+r50Il4u1wFPwEBrnAPu6LOooVE8mDehGfWUo0v41SaxcOeb9ijtt0CUu
dzAfjmY5OTHYyETp88nXBG5zHlO3KfNDcV2K2YhCbqujqUvq92yNbS5Ar9Rd9tYesl2C7zDKWcdK
/qimPL14wROdwU9ZE8P3cvfXEGtjf2zRbuSXdg19P0cbcJda2JTFheUPNo0VJN4q4ocDhFCTisXC
tstU7LiNfdTZ97+7Y/KG/7u7hi+mUQBU1SjtBE4ngWSW2Y0DYpl5MxGcc3o0jcwx1zQiZpt65rh4
t61H1c2eE0pMzdOI5TwB+W6f2//32Dvbs+nofsQwVzKSYSpQJ74pTGduVFtqIUoWJ5xG/lAmdtk+
wK3ho28rQfh6yYvdv3VehqtcXDJWoron2qJDM5teyFt6X5m75Yv9eIHWuDpQ+VMj/Mp7FozrL9+U
/uRkeB6S5r5tUo4JTm7+g+oF5oFUqswfHL9Kk1J1JWJ10v5VeLF2pjmhQHHJZsrwUEiRLJQE6IDf
vXhIEibwwrdvX9bjL78g8iOEpzhOMTk87hwymdkqmiynHhx7j/fJtNLCypoxqJe2tuuhzcCPKX/Z
NfdSBRV95VqaOXnvY0YLL53h46Tsi3nXFLkdiaSahvt0s650sqYsemF3XBTADwCrc6DV9KZcVZlK
51cLTlx/ZLVobBMGC7ikqhPd4QjBsR1ycI8xsIUdZTpEGh7/33/j4hEUdLkHmeZ7aBEpwHpdeLFR
3HHXh8ktDxCm32TkQ/EwzNUIQeP+vpn/lVkUuUDlcQbAvJnUaLwgExaHkiMknVxBw7xWB2t6oJ1/
4KN/8AReVwzJyySkONnwWYoSXQb8licjCW0IlIfijpAQLNlpiVpdL2JFnzxa06X4z1VcmIAAfMPK
UTz7CPkWA9uE1gbsLzUHNl6pg/UNcjGP8t3yEF8efTj3mlRWqVoQwny1Z9fA8C3sBLK8nXIFqRO4
aMwSpjnQ1kgv4PMNTWYgac9AIOuECLRWRdfDKrxLnBrBaafl5HqUBwl2IAFuHOZzlMVSj6IYFGpd
o+aIcVWEizV/FrTYsk5zflzeBNe1Dvg/hHr/L7wvzcW6M/mI72CyJr5RBwbbVif9wtme1TTimBLg
arWuC2X5rreTwru4ecoNI+1JBXeEPeAKYOoIiSqp+tnxyTm1eCbheF4BOTGBqVP52JWN9bod97qB
9fdIDDFetLZDhAF7MTjhXXFvR6023zI9WnYV+yVt/Y0R5s4LoqFWWk5in4hCACvw7wXWMra/XSi/
g6fDCnUAHfThIq1YXbvLba7YxyATW19R2yvHaSWxy7rjpuadzLegCtcRE8E4vtMZ0MkbuTJc32UT
1OWg8ZZ8Q7fCraxlCNg8wmJQrQI0z1RbInnQbsc4clHHC3WRkZ/XsgpvrA8sx4F/31NTKXs7/zU2
TYYixHgDD2WyPQsBs2gJ3vkuwW/H//pf+itHuzE+N+7oxfmMoz5FWPBpO5ZQR/zzdPzaqPaQhWmB
PL2HfXQHA3CgiKHq4YiI3V4G+DMvIFW2QBy4CXPS13WvMpNkR5cU7sEYdilKItG4IrcMAkaCLPFO
urLk0Qv/khU7omwPgd4aZ1dNAVmqlHtCoLgpUysb8JIRboLtzZFJAL8hkHIfV5lY3cnt+UbcV2sA
MiMR99vlNjP7Z0QDkK+JHBstjtA5UwHgI+Rsjd8BAy1GJkPCtSROdxE44EL7IEwPA6AqxZfM9m7f
piMEhCu/ZEBA0llBJyitvfwRuYnMP8ev68XEJHSKL/P/B03ma6Vp/ZAbLgPgbVdXea1nRf7CAIiH
695TuXmce9q1uuIktIMsEM07LzwBHJFxJCxZc4a6rvle5xwBQfzeqfsGtUH72AJw02n9jHd/vDK1
s5G+le5Oi2mtKBNqTFv8sHztpOguToIeBhUMiiT/6uDQ3Su0AHGjYPXKfpLoxWyumrbz1WBGw6jZ
yutVRbF2yHQm5o/EpFGqlFqMvB5FvuNpXUoDUkdNgX56UTXvD0rxkHL1l5qKuXQ8j8S/r+/XcNFc
KDUW8lR5avTfhE4mrzlFBJu+PUGDNfAfXu0CvobNXrI+diNOINsrB27RZ5IsXaIyUf0fKhAZO0Ob
gK4KafzU/9DRRpgIht0wPEtRklAjD7Vt7eqMUFJxKdniNnWPTwuEdlmUilQG5ytURUiFOpjXetZP
cI6EbMDE8aG3uIulFpG+0/45zIshlHV8SHHcNliFllXLJnqynpFkM+COA7R0AzCzU2HtajsUD/H8
skWhl+q1vsxDOVWLcAjwPckznCGqbp1kLry/r8FRC6KOZmI7j71QPlpHlplFizRbiZk+yaMB8fuE
lnIcmDQ/Qs0/i9cNnvKV8Kpq7AB5w5hQfsu0bNxXZUmP7sDNY7LaOk+kwmTMPiUbapOGTtIofmBO
REydSSbsJUE8jLspqYzrUxlGJtgzzKxE4EDXLW6E++UCkpgNCfb8E0GgwgeacSDtz6cyCmLPJvdb
981Xl7bQR9soDWnuFgna2aNEtA4FAehKmIC5W2oEgdNMEurusgelhqN7RD32FrVUudP6KHkHzBvM
4w0haTS2Qywx9CI/3Ajz4KPiif83dNlMzDe2MmmRZRc3NGrv+sBM6KAad1dKoXNxMznYob4dxxch
dHjX5Z/JRDm4/NNdaEDyUz1ekSJ208pb/oOnzBIOamWeYhRjj3hpVdz7/uLVO5Usx9/z38gFR9TY
KsOvEFHOtPV8AtspuVS5npJS0n8iEup9VeVoK5Z3PbI8EDWwchf7vtHEQTbN0fpAwXRzZ4+68SYj
2EW2AuanwstRxU/10xOUIB75yFd3bsvaZRxB8aUWyIFejychppG0geB/VyS0CxcB4TQgyWQvzxJ6
x82DSxaaEDIxoPgnf8W3O5zn+skrUb6sLKbTcZYTOUA8I88q1WhaO8EZxLIc8y0SoVtDFn8qmVcC
aSXZYbwvJ2Yt+Mn7Ijft5g8r0uRuOBObOa4p12z+VciiUrhCBlUkmsBi8TNOqxUhD4/3rUTaes2k
FaTO1CXr+uM4MOcp8oYajgRdRZEcijd/+ZYKC+K9u3Lr1PY8qtRnmsvPqoJQi5etjH8B2BEAcIjT
ZGsyKStfwAkgmpXE4KlU8wK6VIeA4eViY2dD9Z3NRmGeELYHs3sG1LLXdbeAMtwPtBDUiZ2zgNBI
2x8GX8xktszFZJchoxJ4Cayk8kgauH1hNORZLLzN3ZKlMa1O4H6QgBlGh/ilruX1XxQrTF3LJDrP
BKlpCEgy4OYIbERGPY5xRsBmWoDBv5TbIJJdU6OfgtgtaBYAjZSzaY00NelOuL/equKVtCxMexKD
EJr9aoWIo02V6CJIixlNUH+f3Pa5zvG7lDqiWkF371zU2xRMC80ms4sP7VkswkUPpmNyFAtJSHWW
xIDRlknpyuwezvkZkEy3XECYSQi3CJGfZWT//qanu/9uDCHfpgvY6nRwLY6YOioXXigBowQU/fKQ
hA8CsMN5JN4DLZ0qja0ZEbyosyfm+aaQR7McMgGnLMIFf0gdl5Duewwtw0jgBFMn9Aa5VsKcqdSu
Z2k+i3SMNdbc2gFydKSrcaWJUJWqO2ygIwejSmJ7UbTpGM5XMBvTbor0rxhvVr2S9GYNJLr2KxlF
f+4cXkr5k7e7LEOl5h6v1FZ7XgGju563WOCjFdkcDDfPUGYY1WFmxOX835QoKBBR7YagvBMl2PYK
qD76bGqXFlNnWKteyGKM3Q2rglrmPY0Jx11Q6KfhRle1+hlmWLCNyG729LvtzJMSaGU+dowJfugV
9rLKtdVLIDAszbXmOjONmsCvRwXdxHQ7Sd3kU/NC8aL6HHXs+3R4P9j+wYTf7ECIW98jaa01xSN4
9sXreMKwhZE/v3J8/9BkVuskVeRqCvyWXeR7vf7t1UNc5iFOhWe+KN4JoOmiX1lmoryJ42TAhQv1
lNIkkj1jHnXUw/bsNpxFQFuraNNvH7Uo5HSJ0HACA0j+ksEe+WYPrf92Uv9dFgCnIJGwAGl/c8iF
KjrPaL8A4RF8YQjEYhW+pVhd9bEqJ9frsuiq7D26gECelVoVMxx9nHF76E6R8DuTh7wIR2pa1eVk
sgyQ9AnXKAeS/M07/+IfNc35aLvpCOjn4F2L/Khre2qN4kX5er/7ajOq/3XA9ji/FoVc8YDHLCJc
2lLEP3tpO2TFuURH+BZObeoHhIanEs/jvQeOJKwTs4dS2mdTunHt74hFHDjr6A94fR+ANjQuOI24
r3GqSPGCOiWNG7RuiCe6yXjPP2pu9xK5K2cTcYkldZFCvzmpNlvNk+KhG/6biNn4kLV1jPMWJzwS
9rBM8AktQISmkRV3NLKbhpqKxKkajHKI4pbmDUD/UuEdsqbk941ZUiPoxC7K3vIM8g5t1niMndMh
5Jgy6zQ/trgioq3zNclk6xKtrATHQqez/HShkQafUxOQhfP3y1Ma8fsWW4wU2aY248BeShh0hIzW
yNXMF6pgl9DXpU7+B2mtoWXCKti0QzbP5W7Eak/zSlKcjpWI6wORuzugircGulpjHL9pFIavE/I1
aEjVwvuwlKhUm6omWxMbEq86wQNw58bURB+4BrRk8SrdsoLHtO7k2BI2BLegoYDSKiIR5W0PGNzT
PxeEJ+ueGtIh5zqGwU/WvmRl1wtOL7jHJh4ss0NyYsJo36QuJmIwoBNWchEDIAWB9sJ0BObUKPu8
lwMJVOjdOZ/0ZJhzh26AGoYb1Gj2X7PRC9eQCYMLk9J0KU0fqNKjwOSK41pogeLnFvmcEuTGRFMq
hl2Fslz7UbqjyAdi8nlcW+yroXuPu3lG+jnrrVle1I2DqagzoFFitmT+1+EB9RDSXa8QIajXoWKm
H5OvyOzJkagVj1kEuEsVc5CbhXfSBfyI8EqmpNcnGgvWBIyqMumXy8dvkP0JhTvobAEGfBvztNy6
tCjR0URKyu0cIqoo5oPHsI7lKEsoNA8PDpSNm41BbXZlnzI9BgJyfpYZcMfG2y9VAzrVftPENZz/
feSDbV6TYyGGd+1uzewvgzy1vo2RXsB82Jn3Ye0X0WXepmtuOAZtv3ZUJJoE3yWNaJgMkO2Y6jrq
LUR5xXPbSO565rMFwCPBucuQF8zNy0GRxI/rmsqlxn9ikTATDhq3Ob456fsfqB8eETDWodoPqT4f
AC7GrXnWNhZAsRzAm90aQ++oF70bhVV5WH9ci1B0w2003q6WMiNBRUk3lUHPoajqcZbd27TsBOrj
oQASKrwHmjUCRg5GrIuvrVbJhgdAYsH9r2t1mTcebJ8kar4vamJ6B/v2gUSIUWE53FtLH24WC9Vy
8d/MLECUszDAkZRq5k3AadnXtfLD89spy5njRX5v9qP7AIWdDzibZrpOXkYb0568THaKmqPDmGN7
TW1fD7RcGaK+Lm5q5GcKFhRhmxYUFbGRAO/snPxKQEWlpCSXOSJWxZlHjkiP+PaKp0PTDIPAuKW/
im9uzznfKufMZ5J09LZspBwcf4J5l7XHotTtqO6aamyvemyOxN2rIYul+pnZ+WAk6LBWkYOxcjtA
bYSfATCvavCqcPaRvLmsJ55ynehXGQg4zYBwaSGgOHw7AYmzyniz4XAyukW3x4WvcdH+H9dkNKue
UNwRuZI7/JpnlOvM4LU96sQ7RvpIo5crcLR2HVhSghVeKv1ub8xrQBR1Zg/4iy9dSarNIsKUjIh5
rwsLQuWr8mfzPS5kVtFvBlm/U1sgMNAMS1iYXoM5DVOwI7Utie5O/00AhO+HgzttsRb7Z5YasYCZ
Y/US1gqSzLwk4MUng3EifSxRMMp/EbwBX0nDWZvrBv6OScsuNpVqnLMZzLqJZI5fqfi8j6fmFgU+
lyFYEbClEYK0o1GGxBjH33NEPjO6lf4eW47P0BdXoU8qJm+7HoefrVZRAJMIAvCA8qDsCrDFV68n
5C1GQtdP3HXDchnGGFDokyCw9WWue2q2leAlRRJRMf2bTGRm07o3zWLxtVSJJJz9BvN57HG636h3
uTJT9Yg97X3VQTUhmtVq2piwC4+H03I017Zws5WW072uk+o0jJfs4CgcpACtaKznmLloUykHfoQU
roF1CDalnc+KcfNyAbMWjUYO8f7+qB41CmdouT5BHuOmcmjeKNiLav3//tVIzDNxEQXqfXSCgEsO
7LR8ZAJ9gmCCiaJuIlpmIA9gWfMLLfR0cirPBSQm7yv4iU5/cnMPhNRXWwQSK8YdIVqz6++ABjTj
ENopFa5SJkERzB1RwTqcrH1e06jISju/EigbtTrYzZFJ/I1mIYK29FjRQMptAab02jRcxEAk08T1
goTjx7Ncnz2wUDKky1w44oVir9MXPJzVe0kzstUDgJHEvyvzSOn8mVp3EHxAIkwj3dzDXUnje09D
lYlmlR3KS5HXmfSedAwpgv0tchyjJSUzjzVwqxx83UnsNOyaGZOpxNMe6ncabrOuMtk+iH8uTPnQ
f62WBc2/j9VVxhwaVZEbZTLUdT/RoTit53vR4gbbzMxt31pRhBCHKGCkJla3wVL9gVLyfhxTokjR
LxsfzYTFr5G3AD0qdOJaLiRnNZhdtt4FFNKi7+hFPEL1a/jQFpxNY3wYkZiJuJT+NGenVS/IIAk8
XgOvTjeFe1M2TU4hjuehYW0bf4MSS3nfC58kO5dioZMKnVcL/mH1QSo7YYuDVOwk2UGihIgqVkJ7
yn0s+o8ilzuMoR8wnKbqtCP82PapQKcg1AtOm9t+3TgNz10YMg0phDAFjotUrk1yUH9AGMvoyk8K
Hdg9yWoIvU68wG7BE/VViZI+QC7ROHjDbXKAmtka/zcwX/N4ZMWfsMqLt77g/9o/60M1157qR/1t
wAGXnbu3YJGt+YojfQuPQTLXYBxjy3gcvXTtmQOwrqY40+NjBbz6aN79bdCMpzPN3cDj0UVJ7/rp
bZ6s22Ht/IRxkAw4UbYVYFGXeshiG+xmZ0tvP3+c3+SlErBFXwGoAetTTskzpJQgpQuzI8kM5XPw
UxZPhUruWyCD+f6fEdpoE/w8P3rre2VJeXxuIfXpFVrJ/4eEtPgjGMRvFpnGsDsB4XKm81P8Rv3S
qb2WRvzSBkhyuRf70kJp2pulg0a0ywitOwoAjiAWnEOaUpvFqmuH/HJFP7zKBjIyR+cuuVMkYS3W
DjcqYrVJ3FJkImzb3txkgthQdneZquJqn/1pCdW0xT1ZQLOvOIvixYzD4rDrd6Oc+/+Q8R+C1Dd6
edHnUytZc96n5h/DkONxgxaUmQ1m7u1H4nzekLUlHEJ2HbENpSHd8x8IWdQMnVm9npJ4x82h7uAu
Y1bCi3cv8vZv72UasC07dhyk3kcxByVpm822p2OI71e1/KBi7JY3XlW4EE3Uy37fUzU1NRQOYgKx
Gll9vDnh3ZO3F32UNsRs9cPQBvSQVlEQherkgHKzGvX7NGvdeHrNp+7SA+Qx9sW+xlFSChJwof6c
DqoqQUMAgTTviCezBIVcbrZsxNgYN9kL764RYqxbSSKaLLtX6X8JSy+XhE8aBdmgCcDBvBDeAYi/
h0p77tupcj+7l1bxs8U2oNLyEgCK2U2uGWWjnyRayya/INUGZDRaLWDNumNbXjsWx7XATOLlvohs
6Mj+EbbWzfJhLAvgZurNIet4znMwYSNLV4wImFJz3z9VuCwC+TY+4BmJOrTZ84qoQZGn6YOeZ/j+
cUHyVYc2+n7VREINjSC270ViLmepIeD2z+f7Xso/u53sfTmnGACYZnzFAOM2ZOf0fTRvwFMNOHFs
dPlH5dMYOMc4RaNBXgTjBYadLCphYoWj+mlPouSJumm/xRXifehlJVwY8Yz2wNUigS1W/IBxpOtY
Xg8Q2zWoapjEkA/Ghy63si6pKS6zbrByTOsNxs/gthMdeWKpYTbZCthEkwHXg3dioshNZPR8I7Gi
/PdJWhjbJM/HTyeWSxMuHEqrroiX9u823noZO2tfIRBtApLMsWNhqefC3tJU0Wm1J/Beh0xHY3Qr
has88YcKA24fJUEktg8GP+IYFkE49dAdDT35LxGuzUigsSsyt4qEK5JR8DRMPJcfz9CsgJpaCahM
DZHi6ejjPxmTrPAYkv2JYHAl8pQUTxBoYMpPmYBR7eQR44wXx9MFqRfOox+YSR6EtH6+0dW/038x
iwD6Muhx0E1DJ580evtT9EB1+MmbOefTnI79G2NZJ6e1Zt0OCgEEtJYdnVtnzc0NbN0wQgNjW6Cu
XppaodDX/MiClZPNcLF6q9z6Wd9OlK7qI8qYFjfpqAHtzvJTHPFkzUQCbYALSMU+JB43VCOHBTJD
fs74+AM4D3Wg+eMTFnmFHcJqGFr00Zy6t6l07vhT2jVcgRN8K9a+rIstphWHHT7Hftf5WoeucFAu
JGdOFYVaV9DdzpF3sWDTPePWbcnHCXZpyv5cCSh4Lx+3iSE08eb8t1lyUdWZQhEzf92EsvOAFIfM
u6R+kK4d9E6vt85lVBjc7L7F7ymOIxpl57ndB3BKoLQu1xG20HXB+qtwpcwwtxsn5O598XM5G51s
+7teQyqJM1RIdfNOLOnKFlmFaXaCfRX6SfFC9zfAVCu4t9o2I862j6YksNrrRKST+mMaI1rwLgx2
CTdrVqBsAfdl4YEUqZBQR71q1NcdkOPJ3AypoLpRNAEoU1HEGnH41GCuFMB4NLGOTvIeazPmtsxh
2tDZXI9euLnwal1a0OmPqJKhulueDbxUDmJ/Ke6Iige6DinmVnioypa8pmf/yLYXv2+knAhMTEFN
UcnXgWOLx4yQyjMfZ4lH2pRLLhcWn6hT0hoz8KPreftS+pSqwrP/ehBFFLJj8gKd3eZQf0VvbdQr
Boqd+PJiBiDuKNDex+9mwj3s492kQ//Z84K0Idh+BYmvp+zfquKxgeo/YH7zvDmeQZvXaeA9u6mN
rKYmca1tr3ZJIRGodq6d4f7QU8GcXnA/MKLVLk0WB7COyHnRjQlsndKXZTKyHOHC8uQ6K3Dky3jI
fdEJvf+cMgIY226yJoovtSNLvZsEHidKELUD7BrGkpguRqb53k1lBbBOCgIC7kS54HrysJ5VHnJw
fdSy2mEV5uGGkGvcWZYjiKM7g6X8hrpVJ4LRJIAQlRe17wWCalT42IzcUR7gnrR/irmGQN0XHdFI
YucZODDt1Cva0iZ2FK7UU3QvUEUPZp6Qujdu8FxsX2G8jwRoGUiRUvOl0yzNxgQHuMuA1BDZbHLX
kfuX4BZMC26YZp+3mQaAbjh2QyYbapN2OS28qn6xB5QQzgpj1jnkblgbjQOXYXX0wxza/vlT6dd4
iPNdqBc9TYH+gjSC0DgruVMVWI/ST6LuBjfSmLtFXwnvO8ooKaBmh+WJpg+b6t2wbY0ZzmDEwNgE
e4/jRYPXyyFs/2K7JiX8T0SxMu6o/wj2tIzoTnelURLy5xhIefNT0t9klH+8d6R/fLwl4SyGIYiY
Iedzh/bD4fF/mSr4w4+LUWBeA+Huhp1n7xvHwNRe2jy7tx4xPwpjbVCPDXjo6vQVw2nRS5LJ2ics
Vazyh+N8jXIhDRq0ZkwstxFjOHrRo2bcRSk+uZ1ajYpal0865GMJCyZjbnsKEkgxQuR+IKWFfjBE
Fx4zA3gTJZJPwwdqeBqOir61mMe7Ct1QmhyUNJAE2dMkkWqjG4XhVe1lKAJhQBE+u46f81AvaVkM
3Yv5mm8pSN9LVwmxlAOAETlZ1aUC/ENk8TOBDNrbujnarA+KWveooWynfmO3BEh1MTn/uofVuArT
opC8KJ9QU1bmdOCr4M+YUSrUlfDVV9bRAxKl+57YYmQ2jFZ0t9Cam4Lnt1YymTsRh7voNVdSz+YX
ug3oLn3C7LI+k9YdfZQo0C7MTgH1mQEBenW4AsOmQEq43jFywRkheX5lg26iUryNPfO33Lc34Ce1
hAV1wJUWaXF+NXkKRPORBaJxX0t7AWzh3k4heIUatyfdCFaKmFsCF1wW5U5j41ehYMNoOXRy0Q/N
Uh7hlBqlYkQalNt2rSwOnFSaQvSHBngJq8bSohiWQofBOq579vP38VnMkiu+C21IKFryvgvh5TBG
L+4c5Zsu/BV+Sa71F2ja2lGU4aDtntPR1IfAsmXoGtlhfp3heikDxpdjx1MucUtzzCuyPL0DTHtH
/VMSiBmvxDfnRqY374aBJFmrVGOeaJWfiTwXDlRvVR+/So5kKjVltDel7UpRoF+cP2UUTsdGCCtC
8pboXn9AUmelyOLIP8RDzZpCkBWdvQQUxcAlXgsQRQ7HoRt9j3UZcv6aEQ8qBeVPqqnHICkE8EaL
91lpTWYQuY1bSWCMl0Kz0omvHahoB/OR8AYYQyIegDcunXcUtO7L5bBuziyrrHKBNVleP0rpTUWw
jJ5cC6u5EVpCK8NMpwsJzX4sVJXh5uZW9qCvjyxYGpllSomPArEjBYJ59kz7nnAH3WWYZgC2bySO
R6LjW2q0L0YBc3oa2lXa01wa8vOn+M96J6x0zEGSOCeB25V+VMgIyXHjZFaZHj0w79KIkz1UBFsV
ZSHIEqAWzQJSY6l3Tfy2K9oWL0gdsMbNgED2orve66VdsfahaR1T+RJ8BYcTiouShlYyxIEOusQP
BpkLKOLknPQ6547MpINLMZfSmwlF9NyoyNfjMfrHQOR2H83xd248YVs+am3yExZj9RyK4nr7vZww
sw48yQb643fJsmV7sCg1oXQBLAQRG8KWfZ9ioNdBicM5JP126LYHrayMmr7J0qe9CM04hPfVn606
bcmu15+ac9xmNEZhRQyFIlS9DhS7DqqFiFY4h3laaZhzD5RElZcA1tB/55lLYXDnzANIqIbzzbQd
VhdKxDIREqyYUFT4mloFU/ad5P4AxOzh0Bnl8KWDjKuw3VWzZoPUaYwwMFWW1hLfy2jx7HS7dMhI
JxGUE3rwdOCe+DUrqoz9O11ECB6FIBBg3ZLBzzC36toyeUql7ULyfyFlmf7T1owl6sdm77XhcrXC
hgeqdJYu98N0JXW3LCfRwotwNJlq3M9KFSuNelftEN5t6B3rPxYAoUqOoOG/gtMbnF+FnireMo5g
Y2PXR7lVhsW6YstG2m7Va5j+VIDYpbYlvQg2BzuhnWSROQn+JaO6WPkuNymj5PlD9o5lPpux2XOM
4cGJD3NgVBhgxQ9yXYFSLUEW1KH1gbK4q0nnSLNgcA6ZB8gGw/OZXB2kbzlSj8trmfaUSunP1UIH
SPMolBs/O2D7jaJ+1fpqvcCB5mocSMhzYZo2xfuE8sTUB38dGQtilyAasXceJAPiK05TmLeAP+S+
SQwhprAGaVkxrHoCJF7FEsBHn7PRCGz/GUWAAlOsSU5VfiwnEk2WiMIf2AERLne7BXQfQ7DGG9l1
mpikVkHv+AOk4RuWUoZfGGE6oHjrEAgbEN9V1C8jN6FCkM/wVaJ47Pgv3iwafH1PKa+GxBuuYT+H
fwdcSJ1JO5xAowe8FBSL9hPJpN91bjTYl8SFyZ4M70kFKPdQ19wUTMYXVaaiG8r64sbzMIUOSFhY
lRoGwehgYZNQ2rEJ3tHjhC4WZoBW2Y1eYBYYWikn6rZa9DAENdWssE5W76hI0p4YppUUo6wRGaHi
VQKnQo3CauGml8b6Hq9esBvD8B7JUQ/29JeEbmzVXbq8MOCLyjxw2mMa2136ZaEY4a5H0iiXsKWr
mAsBcoCc1Pai9Hnjz0st3bbiV/K/nVL+5ww3NlUNnFdOcWZmH9Hfo6vE7XohEI4jfLqETxAlCkzc
4U2O9LeNd/2DvQwV0hwfGGJ5r8TOh0QRqsFWLsGpehhjiGbsfSDuEQi7ARscJPSNSzV3Ydfvr5B7
h8poP2CRRuU5DKLOuGgPxoubH+lQIpoygVo6GQhTLotbN14BQzz+x/wi/Qg3QosAVQGYArG4qeXM
bSkc9lr3hqvzRvJRUd8Nng47Okm1ZYaWKJjRvvnK0zYnmPA3CvHx34vzl1KxFZo/atycR/22QGdJ
NV/fpNtetRk7ueUc/kQu/g6d3N8caJCrmlyDM06xMea6J1kcVEeQAx01bQoVQXsOUkMYbQvsHxEx
jOSF6FZP34eXeLIFmMlRc0fVEAsssNr3VKYTgFwjtktzg5GjQvIvCuNdliH7eg/WnmkbLpf/peJl
ZMNxbFrR1ZZZtWWPsAmEQ8zAOPTLu6cT0qkG+n6VaFmrvLNfq3wrd0jJZ7zue14BfVBTovZrzYH9
Y+7hFmqoh7IUDZ+kndbMEqFbkdYu98d489WD232K4LIBU9SX+4u1+P8gRjHJ8SjkDE6Vkwo6VIoD
gQ6WxS6mmcaox34QZMc83upwz3WZE2tB9WzRZiH0mh5OPTzLQLQWfTixh5baH1og7pgdJ9Ftjg/c
e+4O3mbFEaGcpm837WLA1W9Ps+2tD/qF6B16PVgvY/smnlZVzlXbz4Qzwys4owK57M6+2ZjiCDoT
eWGVTgwaRYymG/ZXzsFXqvWVACAMBgMQKBEZ8C0Jb1PpQShuOyUuQ/0Q5EPpTnvwaPIOxX6W5Xu5
+6g96U+5Erfu3hq4vUWyOLkywN72zsZHZBzu+vxy4QShcUmTTbU2yworCj6NhTltM/0Zu9KzQIQV
obpfm2dMoNa2yhxs/TXiOHLmeOp9oniGdA6IG0HH5mhZcqCLfAhdLy07xWnE7CpwlW+GO8wuHbPf
BXSK3PyCx4sFMbuqlJM9ZIOVZHv2ooVE/LxR5ZZ/pEol5sMZ8lW2TOnExHFrMsmDLjuepfA/Krli
OTraDrveYjqSVq8Z7+UGiPOz7AMxd/iVyvB3W+iecX/6vCGWK4AVqlS3JXpWoHb8uU4TpKVzZVRM
nPoOuBY2Fu8btxFpaP/UoaAI8o8Pms11ys/aWJbzEa1iY9tS+OKR1SUb2qIUIt2j6jyN485Yj1Af
WFdL6HCm/IpJbZogiaBJRyMmvlMEHBpy2ODlFgY+y/GvDVdsLucI1cr+d04bpbSZmzT7c0hycJLc
mBKZocw3Ay1TMntgZCDVzKhn3yXC13X2KgRXW/FD7eGHXIAKJj9vDEu1MOO0I1oIHiu/tfUM/PqW
VwVoo7ku6Qzn/pCdBOpRM5mpb0IGUCVRfsm72M/iok0Xm6q6ZCo7WBuca8l2be3pfsANECQDwwNK
lY1gpKqyYleWLk2zKv5brbNc5V4PEVDaJlhEojJ7R4YnNH/XqtKIIAgpuxMvLtI3sAKgQA1uWNFL
F9hSyrp1b7qtXT8pbPRlZpemrIX/gPp17HEybkMZnGGBq6SR4Kq4dENsEAB3yXRAZHHsKulKfLKY
mGhFFNp5yIjujvPCya2eP74W6e/kNaFwlLJXdgaAsM97IDNvSL6HMaa6l7n2Ab3AcwyemKsOxNuM
JnU83eaxJz8+fto0YU35ixqeC8ELotL2Czn5Mn2G4K1zchKYnj8a/7FHHySgiptvR1ngkRw5uNXb
vdb1tudBMdl8UnxxDJloP4BKdqZE0Kxwx9+mhefHrFYM4rEJeLT6hlJLDru+SeoeVVIoz43JGPHM
6lYQ31UzoQe5rMs+tubCjEutHmKDFzLqYSteCUVjY8MrVI9WchHG5m01eFB+NG30SGDhZyT5rx2S
GxB+xneWzWxkeBu4976mgGOdpekrnfq8lv7Tg1bjyjoL4Mbxr7PNSlScxHe7acOHeLRcEIPY7H7z
Qmn05SUuAFgAFFKxlviymk99euhMxAM6B53FLaiFIjIsrxkm5MZAfmEqlLZmtsyakTv/24jDQ5FG
JuV4RowLo31Bkuc+3MYKB0LtHoe0xHgrcEh1INySLKD2Y4JhwECwjuI0cf5bgSoVmuJ3COxBBdIx
wrAPjKiQ2hQjk+sp3wPUaYuA2F7OBe0urr/+XTNtFiEfOZSJdQLfxsMZXIpDb3prhSBxtUKM9K88
x9si5xfFRxXhQWoufUzpoJbIOerD9JFccFcGKPkXoq8paza3eYjBaC2qVdVz9KElfaLH9ixsoe25
YzoquxOJy3VjkeZHCXfq5bmrYNBVOL0uloU517WwBdh88Hf0K2oLpCwOTHHamjEfjDP8kVxT1AS6
j2bMp2FiIlrb0dp8kMCF8SvhNFLBrEU3z3QRMuxj2XnsL+pjzHXjtjmrn94w43IxVfJqn5HRqSUC
FMHESFTEA7Oo/0sSYDhcYXwOI8lGr14b/YIgTrbESiFJpFUWo/0m9AEI9o7F42iKc5Tz0XkEQ2tr
1RN8jt+aVWYRgjBCrS2gty14IX7wpjDBqcF5hpiIWdxRUsaoc+td9xSMuR0kYut9wsfYU78auJAN
NNWcTbE7y5mpfHb10LN2oNSn4GtTwkRMjr74eY2fR7GAXjKHmqea+MaUbRgXDaylz0kqtpLgJj13
QHoC2u9unLdthUYQk03VPxQSubmitKXS4fZuhJrbypGPR91aVaDiVVZGfCZcLPnB9ZeXTGCqZ5E1
Kal6Pa+6j0VZsEC+PCU8PY/ht6ZBxdjwjAQ21SH3UO+cRkIMDm2k4ScFY4yhcRY1ZKubot59rXDm
G8dysBEmNJ1w+O2CL0AID7xsc2tguxjBGbjKoNZGrszd5zpsgaBLse6qC1fCaIuX19vXvUzK/dPe
ByU5rjz+xpR98IaRjojTzViN/xQJKU//9CpxOm9Abi9jPJ32O/vWYW1f7ruxxeqIRqqEsDSdApqQ
QzNIxaTk2kMuz8GmOiT/vNc1y2/n6NpgM2q6Kzjixt70rCfr6yncm7s0MCVT60teKYBuQoxe/0xl
wlxszofTGkE3aE68A37oEYyLEoZPWtVPQMcVlCr1+8OFflJ87FLKskTwlBGVHPQ38JT91GpL5QBz
QTrCKWV5EkakiaAvTLmY7kni0AzA+xCCOliyFNURAxNZ7cEdieJAeG+pSSUhnwV3Pmkiavpf627k
darh9xXWqdN/hDd++JEFxU/zisJOE328FpFCTs5tlKfINGTf5B4DnFNk6xcOEN1YDhL8AssveCJE
jVUbr86IyWlgsWk9UweaaSPOUvnA/IZSIVROFIKKGxxLM6tBklDE23mc9nqX7ky7zCuq70Z2J2oy
q1hbpBZ6JJMeJs0oqEAejgaQSZaWhwFyT5h9y7KCbJa0SEUoWH/vV3ZknPIvQULHz2oDQooX+UR4
LEMK8xMl8FGy3D58jaLg8EB389Ur48/EeeXfBxP/EBDkf9VYPgYQpH0L0ou3y4FRwlm3X7i+eb0Q
2Gjsm4DqZpA3UAl65wVmMXrxoiWJh1o0YewHFJMs4MEVlBF5GLjEAz5eXNXJm487r5yudTGX9IbC
U/jQ5ElZNBr7hrptjBIDFKHbfB6JAvoOU511c0jaibah/A+Dk2upWzwV5kpGATg2+D8S46HLSn5q
Ws3+vrojbP2Zr9lLShY1pMwc+1Pdm1OasUh8aRXgv4kBChHFTSYOc+eHxXCFDPOnKuydDl2S1yN4
pCWzAWSVFh0k3WToTI/Rqg+61XiPQ2+d43QylMcQltKD/u/WDT25AaBmiiptDj3WaL2beBsTV80q
G4pZxoKZiy425I4/gphrv1Z+1CpA7suPNirUeqiBFfrDPCw3bqsyokMpPYclnxE9qO7tMjETmsIp
kcnvuWbgaeV+kBfLfJPKZz5PLYuo5pO3ZqvckPwILWv69YVI+1vqrrLFcLeUaMHDP/Q2eLZvuJ6p
Y0D0pVee1mFD6Y2QQ5vbQMJx4wTHvIxD7Zx3mSdnK+sn0l+3t3voLEy3+FMeasY++xxHHAsb28yX
Zx4pjFGlCMeCMF2r8IfrHq7bq9dQKiaRf0qx7awbUC2QysB4OZsI1LSKrK2T8zkFx8kSf/I+LGZE
693hOA2qS6FG/OBqoycJOnlTdyPDLeVtY+H4GmX9nNrvp9+kUwJ3eS1Z7yHICZVIEk2uXwnzCkxP
YsX942+xYyF0LfX5VtdYmBVMisjXSKwEyFRQU6DPwCR09IpqPKX1blUlEvskWaOwYDTVG29Ud/ki
SevEvMXYj9IBo9CwANmXXwFxjiauHUqyU+TREjlvdBrS0pWbjM8d0wqTNabL4YxR5yKQLiE9sb63
4jisAO64SIEVmZEiiT9FAS696BdbCZ8myrAmif1iYW7WIk3PFORZ5gyoGAabwG39eYOoSSvSIXtx
v/CFMsVB4VLwzHcQai8I7D/Qj7RfoyZ4wHX9+8Uz/7ur0W2xfi86AF23lfbLIm7o0WYXY4q1iRyc
WwW0yYZRVqbLgP7InCuu1frK230RzpeYybIb9a1c7Wz3IPf+9X1FetRKlwc8+VYzx72Hwgs8g3RX
4iE9Gn1ljwANxMOfvocMCxLupFk/WuBCHR474Ky4XE2Vdky/OT6ww0/54GcKRI9Izx6VKGDNFS26
tUnvK8CgblwIp2LFD0xukbDPUA/rYNjQ8uZYzpJMMzcZa8XEy4ewFVyoAnwDEVDmP6aWzXD8Rl8p
+B+vSB8XiZOXQpHAotZj7t11gLovUfeVXVyPkzMWrPDz/fl7PFzfZICdqxjowdzK63FkvH+gCNAN
dv6EtXjAsKIzdaY69YW6Iu5bW37LV3UFygJF2RC6NqhfjMUqMvAd1bmW3s1MbspdUj820g9P2hRt
g+VlRTuUBoRn2e3qE3Zrkx1gsb/uvDDfz9q87P37X8GrxgApgbzgmz5Ig+jfgt50QBdT17dPt9py
0T50NW73YsKLOqQd9n7kueaQi6qMPT1LBFVD/IZ2lxTgQwVbogVstQ6iBZSKdpWkXjpwPAK6PFVx
L6OVQbHj2Syr3eZVyQERt2JS5fEF6CpyVkX7ZIECRL20e1rfScxHYBBquyVU9QL58PKVmT1eWvd/
iXOKRmTIxl8sQAiHhJ7qiISGWcpksOHbeNj6k4CYcELC7iblVNygPXa/ftkg/JZBP0GAailN2t76
wYt9JQv1ZYcUEBGJVKHK0i790OQ91REhtR+jR7jPlBUTuVTIpSThNjgd9tEQwPj+sOMOlZw7SghE
/E5TJppkZTDcPxSNUIum7ZxawFR8VHxNnkCk0WhJkvMAXzKFu7wqceSXfFQOS/kKED4zLG9Nv6le
eo5mvuiEVdwh2YOhDDsPUFtA73zrZnr/bTQ09KfHIqz8qOaya87frIKCDqwVQLQSqsG2Dvb62QUb
3lq22vcdmJ/k67QTzyVbDOoqc2yCsGB+bluTjeHeKVb9KKg4YY8upTnG+/RkZOnPMzP1iKrWWHKR
aIIRQMXwQ0JQOD1PDXONkvGBzisvFR1xvsYE5RZxDiSu3UtI9MOclEjJ1eeerXvCfR3bwN7hs+fU
M8wW/UObz84gWaU+G2j20z+tASx9IB8PKmMvycvE3P+pCccDaCfBmgQOyIsCRr6Wu7MkgLs/CGY/
YJdl8vbzqaOM15Mf42VD4ugO2kGtecsvGAxcLQBzIi9OXNqRcmog8posiw2E5LzJWSwPLLam9XE7
p1YrmPoeoXocIIDIGrNW4HJYAGSBnusJUJBQeI6YnsycoJTnFNHAgIhd428BMEAJCMWmiqD6imrl
1xZx/EuX4iPdJclbHqAIS2qMcSCwFpxR5XkLcs8wx65ZDm3q7YQBjLhvDrTiY8j2DZO6WEO1r9sR
kbHLslGoYqypyPyngHERAhu6133V4HWmzSzZ0S92JijbNmwW/bt9yn2X4gkiopGydVN+ZAPqFaWf
O3B/40RAV7p4JyQrFza/R2990uigETHPm63peTR3ziGAOD2IHX4/FawbBYlw5B/9p0HJMCILMqOb
xg5qFv9NEzpcO7CCUlLRq1WiZxUr0jMlymSYxw6DrmQVEvi8BDwJnSsHalN9uUH6r/SMAGUp8LZf
ofKFM6kAibBADmhXuRy9hnoJlq5USjxdhV+c0p9/hZuY+zl2kERkPPULHDq6E8g9DDCorpDLYUUe
mPIOeofGkzTeo98JHDxUNQC0L8vb6i3v74zsFHsk9G9W88lPUAC8j7zs1Xjml2V/442BohKUA/d4
lIpd/SGFriHEdDeZpkp+bAArfxmcSZXvmPWnwCBgIuku/kHeMuNw5ml/JwGvlitprhhze3H60+/D
ezYeitJp1q71b/eRiOcURzdfU940Ojzr+fQD/zOQTGPw4uGmDNXz/OBJ6BcLvlPpIcqtEoBGvfY3
mOlFlK2VINzJeLZlzWOvL5NOBwng3UuElpm0aG6WqbuBlq1MT6762Bu2x3vn/sUTWrRvLvlo4YKu
teXp2MbCHwBmI9qelrwKEk++ESGWXnHVn+NLrv9Op+p8fvgsQMSym3miJC36ELXZ7xRWTGdhjvWY
krXAETp+/l3fS6J+bLMblqMzsPOPYaSaRNRZ5RwCJT0m8iUJVDHdjlmjDZ4lK/OvCFXLSOv4M1FW
I5h9LGgqvEESrgbo4mfA0/1YapboFAaxrokJBLpxzkTVvKtaj0nsCadJU+XuaqoKAlO2L37B1+tG
dBijxmqh+SX1U16FUNYuOZHpceT8U468/KRVPE/gIOI6DqB5aD7TOk6hZ3K+CWIi0DD+JhcbyNFw
p4BIasw1QPS7IjzOQSkk3Swgai9kdrAv9joyJ1lvo+uggoui9rW52gBEvfjfHOVbphrKmS68k6Zy
n6wt0gHi6P9AzqfkfS7nqOp1DRmlTK795emhdqcQBX3GljccACShtEWHYSqIfyS/f7k3ifl1drNN
Hg0dzsohIhAysyRLrebTLqCe3jH8HUhheq7GV7hItMuTPUvjhzMNodKTFIQbfGah3M73VEvGk3gX
AJ8NqkMMwCTiZlDfFmrJzQdA/W7PKEjoyrVysFhbdZ2ff36JdK6/aYKurUFww6QiJdTfrG4oTlvR
tv0jYOZWN5DTR92q3PTcu5jswNU+qvKW+CkRllKNUTjfX1vjoJNkfKW7D25x09lWQ2BzgfHxgAqK
UBcAinA8WTc2NQtDsneEKlPcl4p3ZjirALKpM25vwZyk27vdTdl32gKaM1n1gKAQtx+1yq0ObMNh
DvyzMph+ACGSe6lJ/7oOYvxVfDsqMGvERClFW3mw0SHOzmzfdpwylpyHn/2SiJ9Je9qw46NYq/Kw
395oSh1ChnVYxdhkmPvILFWHlhLibl54tw9x08d47YWQZUd04hUMBCVHjVA4bRNIS/CfjdmEGBWl
97LCPc4T0FsH4lXsqrGNGt5SXE6tpamM+Gc8qLOF8n/k2zPVW3khSqy0eqLSMuUAfU6SCkY4yShH
ZVl6kzXMozoyL19uLj3DwCzNc4j52QVwUGNz7L6A/rMFxlf6Evp64nphzX8aostna4EYH/0Pgme1
1vmHOJNr0zUD4gKUl9RgnJjTyNxTQpu3igRtOEmByx6I9NTOnhykDwt3Vb+j+Q/QZOavEU9JpRvz
EWHL9FQHSQD7qC7yTiFRfe88hlzs09jvL5QG7+dA5JqMpG4Xku0U7N0qDycTi8m3PYkL6Nv7OYPn
SBrp0Ij+ZCvcBpFB16NC1uMJ2RZ4Nci5B1aim3sqywzdHum+XYpdLJLf8pxbSt5tThmFzuKB0lCe
sY4cIoY0Po8GVay9sJq4Vo+2FhM7M2SwNLI5TE2nzWwV1AfV2bTpETAxWkOy4ftDr+IkToQdiBCw
3Joe3uxwXRSamwzr5kyU2H7GWBrCL6Wik9PiKT1aC+lKFpbYgKBY3MFeLVYLM2R7NpHpJ7ATgu2h
1OTyIt1w1aUsy8hDLru22fKJ7sxp5RUBXrhr1Yty6CmBw4gqWNO9OpbnlNRLTCjB19+Zcq+3HzFv
uryAuDF7pW7wZnYdahyfZciMONPM7uOAm2JSG5Ou/8PAAwPB+neY5yYgWB9aFAtOtjoW+HtKzlMy
TD1glCDWDOw+D35IxAjvZac/rppLjnLBWzBoJlvYrF3TtkyI+EPE/74//FfFfkE8Qmd6v6Od40b3
WaJu1HbFhOEy+EQXLKhVxyxxxTnTlvnGdqrAbtYGeFOhXa6Xsdqh+QUdS9tMmH7dGf3MkoOzBMIc
KggtJHTn66xBxecE0JURvajx+QLT7XhIkROs7coXvloUup/lwSV0FLiLU6wmxTSXW4kBGzIJ3uoM
0kq7kVamxfD2h3x4ES0GYso8KwoKlPy8Ti5yIwMNlyHv72nv40ECrwdklqQzbGt6yjaOYPq5lOW4
+P6OKcS5UT+Zwg66e9oE1l+GklTXiHZ9Gps4gcadhRcYiZD0GV2krBoOO2zAjsiynZkAVQC9+iyD
l3OQzToSI6OYSbZEIBWRUXk88Tx7C7TRnxy5LQep4D114kYKFgCmsRZ/CxP+cGVOjc0NJssRo5ZA
ynyqxYz+ZMMITO1eXCBsc8QoA/7ybXgz+qLOcsfmwPwmnnQJbz/YigSRYnNk/3G4maBnr3Reu7DP
uD+EJdZyo6XhEaP8TOXABkBcz/TIbQdjaC9perKUO/WuDjtUtfsgBslXa3FRmAhlb03AX04n2PZW
otZWSMMsw8mV5kRrU8QAJP9Ao0X1uhcNitIqSSlB5JbyHv3gIV/PfGDCseOm6Jez6FayANqFUhfC
kizyniIlL9z1emOPWCTUXI+jrWT9r+6z2KWXhj4GFJ+mk982g/AU3js7+0z66BNjc687BSfJwJO+
hCXif1k5q3Aq/43KheCild/mLFcUYBdGfzp32+eJa0pojqSGy0KF25ZIZQLh3ymab+MZXE8ob2Bi
XYbZJvalkt8PALA7YdaowFnkzTC/LWTne655R2LyRzLf1jWrF3vkzVKxY5/IPjv7lKwgKz0Vgn2R
Hxf5G97pgKetiSd6H15N8no5nHdQnORU52p4WKYTH1Q11G6ngmNLsr1txrUL79wBHf5mISBbvINU
KsakFNfviR+Bp1oet2FQv1EJDMYMhvLSclYNG6rf80918igVJx9oK7g0EV9mn3I+Y+HeFdFPnNb2
86gcTDAF28yRged/dIWIruS42IXW+j6NxWhzScO/5rgakOGnSrfUQqVvJVwrp5c6D51H6Tfgrm/2
b2zZ7LcBvs0YsMsRv6WMvwLuHUK7LcTE1Rh90L9FASZdINWdKa9hLNtWHjvJKqBYm8BkwlB5QLfo
Nl7aykMea/A1xg3+FxFARxhqNJ+a+kwwYuP5G7n9LZf5GXEvaJ+v8zgbInSTryQ4BBpx7Nuyu9hS
y8Ll4X6sX4gQNuXXHjG9AMLaCfjekE1/ov4Ft0of7fbyfMqTCkX/7/G/gPRPFsl12tSJNoyXgT3W
nTGvjnCA44xEfqyktEf7Le0/MCBzzaV2I6rB9THUdx9y4lTyeQa/N5HRtustEC9sDIGql3yj7T1e
YbZU2U7Wkv3tdMn4xA458KEjs0ZDERPQMPeG+Cah+78N9CIYDRN8voQOdIvAqO4PYK5Xa4aiKql6
aLSRl+U227GBU6G7qg3JupGWQcKBrKzX3Qs29JADtiwsRnO7iqY6LrJjujMecpWtrtObt1v5WY1V
w8zmV/MlPdRRVLF0BY3JZKSXz4Y0psfVLrt8R+P5KfxKsHePUEc4l/3TwNbnFPV1KlNmx+YQJSM5
Y+WWu2QCKAuyWuPWY9hOeF8QUEP/5p+n0+O+Cczr72+eRDT2wQ1ehwCoAzWs9PcPrC2hg8JpPgGV
oy5oTFJxgPSfFOzJX5eaa4e+tD1bFXJy2ZSHDDvZcCp5DNPrkYJgCwKFzVxSwkaD24jwIFlUEZpT
p1oMM8wEt84/hNts7MYXOWw3eZ0/mqxhwQ9BheKbzECOvAqBU9cTexeIk+JIwHRxA8QwI5F6VK+G
vh4RB/E8lLTcobtiwguaJeTW2GTO505LlEaRd14kYdBbQiqofjMH79lXd0wINVuFmqRFVph94Oro
mam6s7AXz/r+DLOGNlSdTaoKgxHiP/KqKhYJz7eLxpXZB+ERyvw3GTmROwvtPcuSIsvmlRZephng
Gf5PcdvFExWATLLsKxyRJk1C7Lji0mgSfX867SoKQL60zz0wTeZDyc0craqXmTtoSCbIijz61wZj
tYNzvjMzloCoUAHMmuzji2F3aYBViNlxSyVlQg+5bWK5OZ2cZ+x8qUE+vV00LjDwx/f4xr6LqRvC
CYjRM6plrLq/vYVfW6al2kmgglk1ZaT+6Gtf7xotzb92sPcT1+cuDKH6lM6KAsXKOOiE3qTN32q2
8iLwjyFbEY+XNYq06Eiur0RFbw4Qce7KwtlmAg4nD3G3Gv0M8+nvw7Rp2lSURJu3XHeBVME/ua/R
kmU+S4nfTBHOmmxZuUh2oOcLsDA1mSoCZuS4pP2eiilHx1wpaf0nShVB1Mj/cTWCTeBzjFlOxDr5
8YWnK+MGyTBuOII8hMcy4HCY4W6ItMzPB4NoNcxtUr7ilGXxl51vYrx1zrWGFuJCdNHRIOUlS0KB
ARZbeXi+yElAH6nR7Wp66/7rfh8Jrtdjf4qarIejyq4D+Ate29813axeh3xXuhJN4fMaYg39U+yj
LysnYfhhogUiE3ogRWazib50Nk3EVP+wTCUhWqeXwXRlFJSZ/G8h+Hk3mbqrjfZTLDpZDnIDLDZd
DnKr2+COZ/X+Xa2VvAXKy2STJRqE7sScp/DAEdZj0xgovPSlG7LWm4LI635RVtgm4G/rND68cB9G
hW+pXTdPPcE7YmEuinn9aqEPbygKF8FKD0rDwdM0DoN65FehKhMH/MuczA5q9VUxLJBDbV/Rqi3B
0jfvwrV6/IewMhGUgZTq1UdUBLT4Dov9a5ZN/hoxgmxwl6KIJ+YsaOPaRE7OMPod9l5SKKKPt6cX
36bvErIk9RorGticPZFm+j9Kb1DZ3PYPGklQn51cfbl3S4aOv9WfJUZFt9B7mDMdgIAtr1DkP526
Ar2lhzKIrqDLoCbT8jP5mwpMjF4ZNax5i5XN1WigNlWQ2fvRLNmkc28BTE7qlEfrmpofkK0o3h3g
qCLUa1iR1TTjKIcgieel58k4FvfvvjvqS0MWdfpWvKCwRX5Cz2jQ/HpNfTS+RHMFxOKFRjQIzQN8
NHHWDLyfQrJl5g74/yT14Xf5wmtqFLW5NZDr0TXi+vYHu2hz/Ye0JDnpXicxyWQxNZPfXwaU5BDJ
TyTxZo0yWKW7X6Bx8F7XTtU5/RJlWGzG9i9Fu+3uShm7L0aSEZfAYHGXAaRZ5McqUMVdrRGcos3p
GqUbbP8FgFYtK5njf4UDq4UqXKC6cCmifWLgN9WvbiL8ar6LTC4FTr5FupaJmBnP9KK3MoETfWJ3
KfeZxzM+RvxpZi4Q8pgCMbXq7EJDgSiH69tSLERh5SsxhKfbXR3Lww3uKwkKMKjhvWeNJ9disXyM
O2zfdZd91nMCGlDIsHQ8ZzjXkb+SNT/ngkp2Md0S1D1IIOSjdqAzX+gTTIK/oVM3eKYP5jIMr/vF
mBAxwqNr4/0maPMiALcStsFPdyztnG68xMBXcR6G5L7USFkaB7puPcYCIqiE5du5TcTn/qXyxDxB
PH8J9t5ktbYoGwcKcVyExSJ5P4jf0D4huO7f8qoQkzxW8K5417AGoUPocoG5t5jKOLJALBKFPeRr
UAHo4T33Qz2ChYA9w2uWP9gOdbIiNiDwFk856etMVWWrCPVslRflrk8e87q6v0ln5OPnYuo/+GZG
AgKBeXnUQSYnrYBDdfK37gv9omZPox8oA0Vi8cHXmHaxkd3mtAoAMiErMALsaXUce3xHUfqmvwpy
JoFzxWuWWm0YYBNPELBGNCJR9c6VGNGoYf6imYW1alEvDEovLq/zZsL5f0lgeohLEsULx2oEeO/U
r4X9lmmEKj9tRt/arMWKMuV+nYI0+w2n71Cc9DvU3q9rByQPU5gfuRvVxuUlIidbEcnUFSBgBmB2
LmOJKNL+ZVxS+m+5uVOwUk4CZdzpXPHs/iXXuNm6I8p2tuDjDRwCeclFKEFYPqy2rA1L3V7GUwFq
zMPsDssXC+nz5HJAgKQX/ep9VJnbyoVtxAnh7ohY9p5MLpOhMJ8586LWv5lacL6iIDihRWYmYrRF
tmu57TP1DchQIOe2GSc66RP0g4nlCzQhu0kdMjBmFXWN44bIOTGGW6mDX5y3H/EF/P8Vsg4PMmeX
85gaNvRLKBoXyFb/XgXrmA6QQJ4C9v9ZJG5Ifq+zAezXJvLmmk9jCW0JIZRysbx9JynyUPZLT52p
GFD/sEs6URDX3CGpCg5OclHK3TfZlHmpMWRDMfEA2tT7lwfg4CUxIZ/UgooRW6KqQVRYDyVYtMiQ
5KwHzucMHiEEsvYNG+SDCwrC/TU2OM1AzOY2uPbZEzmca+LuETQGVO77e2pvA4Zm8cYgW8rzR5hv
j3WHSiN7wEdYXN14oy39VYa1EgvzAnxND3+dXVNY9JJZQTHfi/kz1zdbJ7z6i+8JsV7HPD8PhZM8
NYiadZQsSZnrqxVe5pfdqXcZjG+epckYciNhlMN8kGizd1YPl/hkbbHsZYxvxMrItEYwzE3I3lrW
gfCpbR+8PnTpM1rxzwDUZCqRPU8utKgWJLbmq/GUtka5OczvmkMKS57jaClskCdOJYNuBhA8DX+a
DzIg4+CC2p8XIqZ5kBUH6Kx/rGyQbzKnLO+sffSr/YVAtmIe6ip+WLi6TpBebV4QB6cZD79mnRo3
3HbUys1LvC6ktytjxxEdZ5YlziqgambthGP5o0m3jKXowgrRtfs3tCV+2Pr2Rg8qteAWhTmBnqG/
2mq4r3rAldkAHf2w9PsIyChV5u0+XJ9b7n8Mb+xK1xUmhqEoppsxL1W+CDTVA2ki+f+EDmNAR2fe
KM9Fu87eHznXIK9C0BzbHeKGlzPXQw1Ob7iIFPPjyhBBlcI+dt7uCOPgZun+UuZrAjqRCzhv1cTF
R5HyXQfFIPnmD0Pdqs9KJ5d20CZUTXJEc/JXXF5iD0trWi1TrEi5VmZAjE2zcZKoq5e3N13iEbPs
uZCP+QvSUWINu9XyeYl2JyU1rbFxuotepj9VYX8vxw3YnIyh9Ary7YTCH/ISD5MAu5cQKHxl1T6u
/3luUExDplkeux5KlHPR19UZ7/hPpNCq4HqiMcOoIQFdmc3e1dmvaVZV+Z4CZ4PXYHI6tTz0zvWg
h1OP163fM3y5WSmP+Oz9Tb+m69+yKyEN79rhnqzuys3XW0o1H6upAnEvN2p/vAZqjP23819eHJ/5
y/SxJb02TX2SeZCL22nRMfzFSerhyPiONrHtFMjM5eI/lydL7J4Z6Fs8x/7/yEQq2MprrAttHVLz
4KvkE5x+f51g8CPIVX0bCW1GQk9iqdjshCCF0v6DUcTpCjF43zjoEzeHBiitNZeEU5fu7iYj/qF5
RQomzL758YEqsbrhcO4DWXI6PHh5ogUQhdfNYsrcVedQmwEIYUrKFSn7I+lvqM5hi9+qBZiCCU8O
fiF7XYaRnvxno47sofaDXVdiHcMUZBSeVrG+CU5j535MUOru1MUVzqNzHvrpDrLsZrzi2qHBailx
M5H+5spjYHuRhN+K0d26dsp8JVsSQfNKnsX8InCZNthb0N0rLuzwtuO2AeA6Fsz03nlI0GCKQdNx
KFv7LRptDAcIThMEXPgSbQ0J362PfHgnM4WOfu7cK8G6X7AGn4eC3UMXLgikzyQ1n7waU04/D4q1
cnya17gqNboeISLoV/VJNxqUaDYY0iJnFyrUeSIK2w04y75pcMsYBbqy43vgoapqL7ERhl2Xc/cK
8QpIcQ1oAZvQVVgv2PXqoBA0hscrqrPaiTot4n+3GX4g1sXHK7aKdMVGbWyipL13Fi0PV0TOplXe
od2iD2FT5kOYLorSDoazySMbNgwIuX7vmy9xvZoRT7vrUkYFvxBlEf5hLJUnzT0J4z1MoHmH2LS7
TQpTQL12qmDYQu0XmvLXuKeHfeqQUzk/Xg9wrSGoMtECPe6wwBWI5a15ibkDv/7MdrMP2t9RBWHl
VXCERBgrCn7sCsg6cohqjRmoxcbUoEe9YPw9aynUxel/1UzSDgsgviBrwEW33cwgyqgKY1eSq731
BFVP/I4mvEVqwWpRKu3ihu+P+4wVrsuj+Ux1qUH0MXYAtkg8S/Vgqa58tCfcaiPH8unR+gjmwrmX
qb7APCdgmD8g5NlVqNwg8ok0K9/qDc/Pw4gNieSUhweIutrcHgeySnfdUOjOtxyu9RHc7sBQzNwG
c/EwnLz5xlUi/5HB3ehqcRG3D20NjNfv/fZ+uT7fgeqG+JRGFeGfeZEjS98ypNwsWV3sLDDXPQM6
XFTwxAdIlcnT/8emL2XXx2T8rzmC3T2U/A/ePnZjfrJXt5cl86RI6qt9dCjyk3xwZkDuEME2/qrw
k9pImu1gzbIxrb4UVfPW2gcgAqsHzaa79dYLtnsbQIpY+CUo3TSmJgvsAEr4v9Z0dEM/OEYT4Ymu
bL19kEOD3Bs0j0vj3u5tatbv4zdFuTotXrebJ8b2tpn6FsDT9CQrED4caLBmXP6QGzX9JH4kbR3t
3ktJ+DSGfL6UR44f/fOBy6EGok7DZrrNgogChZ3ctKsSNulUoSQ5mW5uiChcaBmRxoiOkC/bV4UT
2CI7qgQzXqlfLZJGeZe5cse5If5QYBxgUQlEYaPgZqEP+de0vUABqcBV9nJtgkuPdI0PurjtMi0q
PWjk77F4ciVI9Vz5RMy9AClRbby95+sGFflh5Fg/pQ6RMcW+paXHn0GZWDlE0/jlxiSCksfbbuS1
NOw81zF5VwYnCdxpT4TCXwO3sX9ZC0AJ/ot101q6/AVtpPJVWwAxIkH60tHjaykKkznFI7rYew3W
dyaGTwre4vtqut/wwpf09eEIYLKXUMGvvJbvCBWygGWSIxthXdaisfcqzKcnlDazVI+Ivw5CAbdS
20W6QbCvA8wpFo+8oA+666xmt4YJ/fI85Q+Q3x6Nk6PzjbfDWVtvbii7xkKE1je41yL8gVr/gX9N
y0DEECS5lvv595tdTkkgukRssky/O2/CFSULWTENmFaBhD/TVuy46qD+hWLhrwbky39dI3yXgbgl
qO9HUt2W9YZwkLq+TFurjkhnMNCDnNY0xwt12tYIRKs4dRgurXdQ1HXdpZ9QAkhycMY+K3py8aBR
PL3bMUevlTLTJDB8yV06tLvbf8KLNRILrhFwqmT6nYldyyERZFfqdSbHTM66c0sOIToLLOCZEWUz
OAVoBEs+twxTPFfl/zFzedBT2y3a32KzmgzG1LoZnSlfr8ToQ/ouujnNt4HsrIypyZRR0TpIArfs
AtXtUNAfxwnNWJEL7MpMLkZThADMhI0CExU+Uum2uXmC2OSMltjACuO+m1JAEzPQmCPWBbmTiqZk
0fj5Vyf73vIM4EIMJMD9jRt9DlL6oqJexZbhor6jUblzNfEMwKIiCYWTaX7KxtYKdY0IKMr+W2WE
SfaKa7hW1R6f8lLaKFVEvZAELbwX9zFcVWl9+Sq36AEjGsMoiuPq79TFPptgUH/6FLvxT2AkrZDA
7Yf3r1RNrPtR+nmCq4XbQarZXGqQEYkauq53iv/oThz8HWZ0I68rq/F6zLYaT/P5/M8fKfDPdHs5
7ZoqIsRgrpZPjnvJ2IXQGMFRbMExCitGfDNTw7tG5Ak+6j2pMUqSjSiberkFN7NeMklSMoX2LqLj
p1Bz8y8tIUhIftOnDGYdCJyxIx6MjP2M3Ybpp02ZxgfKoiY9J6+YLI81pvCD9HuufdM6iRXpxmIy
iJCMHGxdAlkxuFifzSEoCSc87Vq8hebqmgdjeeIv5Ni4B6nBoVa35zWCnKdDS0ReDpTwsRYyD4yJ
ls8jq9DWJe+VyOKL5s6/C874Tkvtq7BMF9PmSec9IJiKsp8NYtKRhgBVu8Zo8MDJFkKWx9XMNENh
ssLtdforqfrIWfuBnWuAxxLR9A7o+4a9l04skZOKsyqTZlawHk5I1ihyKBiz7K3L3n+Bo0lyojQh
x2v6m0Mdw392qFEGy4hnZNg5VeCkUoqQtwgrOIkiLDaFzzEiQMEviweOujQXuLh7BivQZkAMIY3Q
X/EMNdgB5LTN3tR+ldC6sMI3zDnuyZDTpJeIClZ8owKi+WpV/Vw3sPhCXL+qbPk4tk91A+hhsAIU
TnRUVUv0KNyfs9k6gePsu5v37GKwbm0cYRHykhvudtwp1Z/yn2zoIueYzcamr1VSdRIXzVmyDom2
FoBlazga8L5yvhOtm1IQm/rOLDJsuiTUBxzhwI+r8PdCDHxor8q3MxMyonzMTE7GAy1uVn+M1g8t
X/ncAVvtRsidEUvp1sn0OiaKZ4tJLsEamEdpoSbsWTaLPydvGtmeMvzavqy9ezrQjciT2d4GzSva
GDDECF2Ya5Ndk7E3/LPWc6JsVkV21Al8t0Uhxr4W9nNpZR+ucG9cyXYp54CAXlU6DHAcdnYnDXD0
5UA9aEkCGVbtRyfAxgzKt1bi0YsLzudsBi1oxwWc5EkwL6UeVs36S92F0GcIHw58NQI7IdjEMYEf
nqrzlrjwXtBDeVUrSHmTjUXa1drlCn1rlaAJ3Nk1oaCaVVnQezPUlwfN8wLaSdK4acoMMO2gFnHo
IiSS53tDpGx5JSDJX9BCC41USJxCMh4t0Kbd9SeRZTGH9xVZ4THQAws60vdZTNOJ6GB7Urng8yGD
Mj37NjiU1kT9uEYxDPHsWNXlnESCTSIDBHRX6rniaeU7FVlqbs+WA5dYqajDliDc51yFL5e9uYLe
bN5FJUhVDlXngnwj/AQL0yUqA8QAcWlXAnuQPcAqJZWvvPeAYg1jV02nNg7bOIU3uLQfuoOiIQtn
Gu9gEJLRpoZ/Y3KuvnKaRuNABBnf5pKzc3K3Uz2MA4DvlkjaQiKX45mmKn0BapuwR7I6zDOiN6Y0
uO+E9jDymaEwd5nD5mdRfDdHjQlgSg2lyY1gyB6/T6RYJzTYrs2YeuSH59oYwIBmxyaIfHXXITBF
F5TkIr0qwlf4TnGq4MyMjCmSG1V9UAqs8e5VykGaLk3fOmngcR4friJhuuLqM+WQvqcAXVC3Kk5G
qesn+b4ybJ0fjYyQXbXSIpMVyWO7zGvJFI2x/bX+o2xbzA+GPcn2trPfY4/fDrYYEe/Pqt+U3ISl
G4S6xor2udm2UCl4512eYB3lYyByzsj/F/JWmuD1ApQjop6yHRpiKo44gA2e1cTzmi3NgZBgODq6
yWY57OovBmm7SataXUg9erfeWaZNNVImgOpv+C59+xsSDOBqyAw03ueP12q3Zd1YurYOqGFVaiaC
r3SU1CJYKn9rg+t9rXeiTAmMdVinRZ6Kg3WX14LIN8nZthNvTdoCjRRBRD+T0SBzhAV0H2ZUatxC
wmzoKdKnNHoLZlhJgT9nu/4Zz0oTGkpJL6dBdN2bnAq63LK7GSzYlJM67ZnHBrjkZEOc2TQ1eMGW
+ZfW78twG2JdMS+6XjBwOg3uguzIKL63AWstkxr/ou+vSnIFWJ6QA/W5MWXurEoCgSs8C5fNiiid
cgo61e1n0n9xYea9inney8EhNTtAKzGX2TP7TJt1wZvk/+TU69ZvSNZ1ffXuy8bGNuLmkFffyMpX
gZvVZ6TL7B8X0wUfmz3MX5CC+lLFTwK74cYmdkxwqBb+YZ4NV9qMAC5sPGmJ67jWXoI+HQ0K3Bc5
IWRk/vzvn4UV2sC+kPivJxLsHGoxZkFv3gsgbMt6Y1+sD1l4ouLFX+2MCMVgRfqIKnzIMBEw/ny3
SugppMQb/O2TO6E3xcs60u4fBkRhArBFK2fnic9IrH9nvHWXMFzTK+FTHOT9tI09Z+6WnVRCICYf
yoT5axVN3oq8aRI6jmMCNE2GHIYPVs/3j+oyEop+R1KyJ0m9bq2iRd+6xvSnjVMnrg4tF2IKhLZu
Y12wThAK+QNYunAjnpeDt3V+9nKqHY3t7GqRlmUDULoipxBZgBjzuqYQ7LF+6Fb6tpkjaVFTBAhQ
dGy11PZqB+xxzcO7sddU/aPPlf3TbuIKcMq2P5HSIgNxdT/XRbkAoyAYLOMtk57B2iuhq6rW9LlG
Rxz1arwrwVOriYz5fEWcuijfP8/v645xWbpAubcTPntCFJoWI1G9JtlYmAWtD+ZIhjvpJAU8fxXv
DE8lRMYJRR3QzcbSyPegP1dZ/f6Cvg8oATGHuW03zN7s/XeUnNrf7W3bocFFpFvuveeDhsrBOXTz
HBWEHJDIxWcqoHLyQClQKBrD7vsdSa/CNDCbSwfQEGMrn5tfwSShQl7sVSa2ZtKQmQanlFWewMLL
mt2pYfptrEAEWDoCeIV0VvgVk2fgR1xxJcJ1C5xP2N1pa1oa9xVMwHgZTF6G9OYTJ7axn5+kouqg
Tv6C05WJ4aQW1gQw/A/eIxDl6cvtWFP3bDhZ4S2hJgBuSHm6Dq5NeK0Wt3c9rR/eMM0dJEwLdrQx
YQkRCeW9s8bs/qQ7zXWy8yBUHwEuBw9idb8nQaDlj5ao3dl6XEVtJ+qFdIP2ILY4mrn9Y23b0TJN
K0i0sPhIREt9Ms1LvGYY10myjbhNp9CriZX2Wh/il7OojU8sfql937B5OiWBthZFmYadVf14nQqA
Ys+EgIPxFqbQwV2spHTD6sJ2CjpdQE/22KEbi04BolwsJeC90IniNJJQrlgST5QIKklk1RUpSa+A
eS327h9it9z1nGRXtq+J7oUXOdF623H74CnDLuWIxi8ARQi/fYx3dICigqQxrsNRFwW+tHoH0H3Q
5PJhgPENKLnN/p/qZwKKomKzp6UaiPD3LztWbc4K6P3+cX+UhcNaRqUyMpNCpqiLqE+3BGuPLH9x
XDS61iyqNwUar1VSDqzOqUGnDeihAPTnzp/eTjMbXU431tOL3wUUsbY76hXUUeeeja2DMn81QSty
kBpb4JXrtnmIreh7Hb1dfnRPPeaOLrCI4jWEZip0Rd4exjPNry/oy2wd7cqtKQvu84+Hw43LHRAv
3QRYq75s94OHt9WJX6mw0vW4cZGXCcqIazTcp0r9wIXor2560V4obn1ZGi0ZZiGIB+hCJInRsSAo
2RegIjl/TgX27x4R/ShHxnQXbaP8fzgFLGSObnCzjoYNMjSHwghWj35awkIngdQGGMAuJuRMAr6D
JGbEFOJx2pAzTnMcJGa7gAlfQqJbdh8V72eBhm0TYXz6ipg+2imyH1xX+2g6y0+5G3SdmH1nJTvp
OfCSo7Gi475+8fZiTiN8LnnIE8Ysk3UDqweMj2eyE0fumiKTSl9beZ5ZLVdiTWxYHw9rXtfYxO9C
qN1L0CqC6Pf4DAHX+Cz6vvLp6V/Y7N2pPbew/OG9xSDVeEuU+NBO3IAO9aad6I1t0fdu0R/uWnlg
KZRXBkGaxWwmn8VyZOrENDxwrmHSBjJmmE24+IxL3wZwBipQ5gzPtXs02GQZ5P6s3K8C/YY1A6/5
hJ+Yx5l2yjxYUR3sx7zQ1KGZ5j55jWK7LKTC3f/fqRa5IBCGqVpg+uSIXzm4cVdnO/4tt+hRI2rH
l5PWE09vsUI746VMCJXEymi9DqRR42MQcS+doc+ZspwQm6Q+qrGYETu7/sD3XNWqOcbsW083LOOt
1qgXGy+k2km51JhxfsUzDZJbBtKwdsbd4krkO2az8OHZ86g4etQBEnTGCNTbpMeYEoiwO1W+YOMP
eekG6c+wIcja0uQc4Dt/ExTzbbtD8FaHVHlcjDXK+yUAjYqrNy5esSv8E/UDugpnMnUHQVUb0hIH
rjxuh935duDa+tfBVOqV+UcMoI5hYPALRnUzB2bKpl/DDdJijN16ESXObkBUEh9oBvxBfMPvyBXR
TEd0+L9djg4haTTv6wrVhpnq6pEhaEXsNSMLIYyZF4ll/NOEgToelcMz/yJRBxJXgj4ZMw2dZfOF
XnD4KbEMhvU/1G6EmmGwKo+FoFNFmZIqQigdzNNiDRkh4cowZRKyw1qEJveX9Fa84yxvc3a5FTFW
34FpE97Z8PwGVJNr9uU9XopeqEEzhpY79NCRPj48ACR4KTEvvYUV+t8+4wxFCMjAc3pzPwes2+QW
16cLhFao3IxD5ukN7qhq9gr+KxwtqTpsnjsCV4sNEk4a1bvlONCKo+SXNkYUA/+BHf6etgQbNU4g
S4MaRU+Y1lX2tIzWPfLXL/dOIQliuYfwMr7jLwhniWcw6+bG9e6/0WTQQuXfY77kP+ryRvnEFS1j
sqy8Fa6rWvFyAlONGlrirT27OJtDTDb3aAgqAyLBVTmy4qbOi9xEslakB+hX9lN+o3Q6KjJx1hQL
SJCiXODS2wA+MchU4Em1Ppf6PoDrMxnpNYXahbxnOBfml/8di4LJ3yAPIkMByNg5PYyuvPtPfarr
mSadOpQF396tP/kXlVrQSoBbKs3wfICENXmf5GrA+zZUT6O3rGt7LGeASML78sWZIFnZkVatbui5
kY3QaTWOHycSyPI+7ftyIL+65YKslsjvc3sfSk9pjQ9JD0khHsi22iYa8LG+z+/10rJ8VQlxpvrF
1yQ1jEMpgLjRFqPc4YbArgr4UiIY/bdbBwGgQrlOhnhQqQI2Tdb5ox1ys/OUY86yGvhZfS5Mv2F2
djXBmfDIOtB6fV2rWRdbIX7SUgpW1Lsj0g/GobAYwvsK8tXlIiADP+LMYiWE0jUPSDAoV7vJ6LSr
3FoCtppOx3d3eDnD0H6dZjwyxBv6dGNmM0WdrIRaaKukWv988vJOy5NiSioBZ8WsVESP6Egw3/zC
Y2VjUxPejoiMc59T6YrELrNUVSCusG5LnQP3nmTrp6S4Z8C5M5URL3ttCa4q3YrCBXlFBRmYNeZH
lb5CQzwEhvt5V92n0H3HuHGBUUg3SE6Ydje6fXls/xrqfSJmT36iCXj6ZRVDQRYiUXmNU6kF8DzZ
BDWy9DXiM+X/KVap9jDnx7gazjQy+CwnvFRFxuzq11YhzJuOcipwuGks1sjzWy/U1z50WFhcaHFq
vg+nQ2gCFkGiGD22yuUC/9IpRFQXUAq2wAhlKCpKj5jMLBsZVrLHM5nR2hxI4Uu8Lx93vwLPdUZ0
5L1GXuTjt8Et59BegRhOjSjq+OVDhCOPpAN5CqOMVOn+prH6i2g878SW4Uf6nvUsJwJjSfLsqG8D
vprSUriCk3icpEYklsXfcO0DPsAyirgWxbl3VQs5ElTv1WxuuMy0Zhb7n8UsNAXkABEV7WCRLi5n
BcgjCE5nyvq7p+zed5kMsKCrvjgHWyfNcQc9NIY8xAV+yv3+w71Jtk4FUrR/8H+r+K9ZqqFfDa1V
ihGAdEIlHqKgaVH+fZt860naTmQMWYyMqaMgMCCEuQhPJPvRcK7eZtmySqTBMQhQh8tvpYFZPvbl
+7VBMQZZr6Msfc7VBZmL2+pvfaO1CXVsh/b/ifNsN/2mamDLnl07wVGdTmznoJjjtDSKPDMO1a1G
sr9UGbImsd5VNxHYpL7WTD9TSSvdQG4EIymCpz98hLGgdy3K4Kr1Auf67UfO/CiewSWqi+yhfWNx
j+WyS7uaQXkmpNRwh+XcG3h4RUDdMZRQkE7wnVVoSjgzynwNe4HgCj5YkSHC/jM4eH9d6x45D/fv
89igG5vepdJOo+W0Mh3yVjmvCkWKTvP+mzejdlPgizetNveQCxfa2j+M42au3JQYoc3QGaOnSij9
Jqy8x0UuS3uJV2sMzFiBh0LMh+XNRjg6RKptz6E5tYPYp1z9CXFjfaU+TFo79dtraMLgTf1sZZTO
jJ7cDwPQIybQjFnWw0JeKSvgsrpZsZOl2/h+XOOEAuD9b4NN5SadfRHBlVfuAmbz7e1iCUkAQrA3
CVItj5GyoAT5ghpj20rIKN/22hSF6MyJtNP297dXJGeLWQ2XlTlelxqGjdwb79ZO5yC3Li8FKXkM
99m1Jbf8ddsBbsBkCCrf7qjP/FuuZh4BMMlEIA6OtUHV37dv6fwaUh6U2oo0Kxd+3B85A05l2ja2
fd5bFmdnRrvd99ScC7GxHmPJjliglvkvCkkjgXYxCRE7vNIPKCJEsve11ouruIu7DlWfMMICULte
5dsMlelyFgmGT9xUW9H/+nI00arx7uca4wRgB1unun1Xauq8zQBUUWh0+KFyNQ4n0zL2tmWRjurI
Hne4ZDWKCAgFVYqAF4kkXMBMwz//w2uemCsqtlEbWP8C9465GUMOMwxs2CuvyDENbbOxKmYbTrhw
n8ZoR97q2VAG/suj0qGWODRy96hpV3naH9BgSxisNaPcvM2c28qsVSBcPs7DH5Zx5sPQtCUo9ADe
SdameLII6UFcWFkTePDrSE5Y5TJ2OUuWMSkETGJC3JoFFjpQXtlhrIBKCNE/dcU9O6JmVPimoyvR
y7ZGs07difCbnRIbN1aCc6jV4ggoXnhzqeQ8b1b3FPMQ9fQHiEfsQKGe+V5QPUqd6cgrrNkUKBFw
DAplUgOmvG9QrjpEa9+Rky3QncnfArXp4qWOhRI+tBrIogA1a45FaTcYuioMG2PIML4kxWhzlNEG
XJEaWOjPU0LQOkhY7huK/h34n365/xH3/FJo7XU8l0J/Z+CckJ8E5wwiyr1aPC06x1vXzXxnI8oc
IE2q4rC2Wxk1fr4LNKFnRlo0F6+cD4d3tBrw9GfB3hgJlw8qC/F0jQ3moX2IWdsIG3B2D7P16QBG
yqrJlMi4wI7CGF0E610czJ73JuURKqFy5Zx389+hfz2K+kie3zaaZZy1UXv0+J/aAah2YBeFq9NI
0CeeIURiyVEE3ZCLse93Ixrf6f/MCY+23VHRhI2ATQt4YwbrzNx19WQv9YQc7mZ4l+iO7YwRABan
V3KeP05RR+BGCYjBfeoPODKdFSLeRk8ZYJpU3sC9OAwQD+1uTTPByx26sUPIhrisNHf3ZVo25hrg
8jw6koi+Iq1bQUhB4lQ+U8YoawlO4aJU+LkBNX1XeZ5QN6J4qzgNfcfWKjJkm57bcIojoPNhVVUf
//uF9cLdWTa8ICI4r903Ez7AN2/cXE7Xy3pQMIb3LwaDIFj2sE92Go4bEZxwDWiNUVxcM/8IstU8
mJBQtkns3bahEiIFnwJ9LANZryQhnfkxS3y5ztXZwT8GhleWw0Cvv8fg3sg4U4Kb4o1KKqXnw4Lz
uaUtLFORHpjzatw5v+QSj7G3t7jW24VgaJuLIb93QjvHUj7yjSfjI6vqDiw6bVG19houJVtlJxtK
/8WK2Vy2esxnFq4CiJhe5/he97E1371xL27Vus8aHABCtweUZwCQrEjWSkTSq5xUxe5e/lNlFAao
DqDTPNxXQ0yx6Q6q9mwLPK679Jch3MsI+6YtV+UXDzR7zJJyOgrkA/LJf8JBrWG84nb6Npue6h8n
fKaxWuXa8Jo8XfGCp6GgSdxfqq9n0nGThjEytDeqCjEZZFqeRuzEjCVs21oAQH+Z527m6radoPwg
WDcRTv0fQ+dvZOwG+rv91fvgqjNG+nz7ZXNCh2HHj5r6dI3kuMKxjVYpfxIkcxXFYIBAGyE67v0s
XCQk6BoKGOw7hbEomF/wVE+I57fG+Iel4biJI2dUqrV2lOUD4Gv1AIwTxaqqO/246hkyxLnE4+Jv
Qg3kOqk3Ah5tHvDU9FhdGR8RTyJn30QXUf10VrbO6PV9UtaJq7EE6nwsL1vAkROwqOnICqGiCdny
prwst8g4BsMOYckbih3XSfaF53hJ8oQ7yra6kQch4P8cP+wj4iaWFH0DXDktel5JCIvxzX7iN6qh
IfVjU2ZzdEHDzP/em4z7TaA8BbxUHGy134YSYbsaX9UHlDc6Orxghd8hN2SaGXtNYshAd3KqCuZz
hlKdwKXMM4sq/soKK/N5PtTB8LJeaf9DLN07y8CuhaLBaupT8Va7LFJ75HLWKa8VXJdff+5AP2Q2
iA+DT7iktPEbP4ktm1ORlwYpTolL/GIKilHHs8Jes8Na1CMZSXYnKO6KcNAkASVrWv05VYciEFdv
QLM9IAtC7T15EVaW2iUagAPBel8g53ey/GozV/zdejZ18my5KQYH9bGphsxkNrPE/UShx0P+pGZ0
0vai5AzbnGdzmQKrqklOMSaEiv4G7Esu3CiiPZquBfPxRaT1ErN5BIrDcGWm1n9bvvS64ZOaMACc
7eQqcCTReOwMrZU8unISXk7W2lMQ3Jd03VrH5YHVzL+x7rOn6SmP1yazMfnY2xCeTqT3E552B+HH
flpwK49giXoJn/OEkc0BD4L04FAKW1TCwgpS+HLymfa1wYsNvQ67BjznMTkfdl5poH59r6CVSnnc
8+nbXs8Z9uFd3G+kItPTRC1kKm/znlS9q7gbd0MYFKQT9w7yzvRQfOxDxzQomFP7rlDQ14eriQfG
VhfsUFFfxewWB6w4uaS7PlWGgtX7U25S49e5mVWkqE7ItkBZMftuITqYJdijQ6cBW0PIOAFo9Z9r
r++o/mzErn3JKY1qxwAeVZ++iKAZz5KMfcyDzYMf1uRSluT/Kx+PSUpS7z4VgDAcVeaVcH812PA2
4xhHOjNwdBGyh+YAoOxVChyIkXIABrKJB6icvPytAQ85cqoIZNCAzosOwLXXkA2O6qbBT6HrXn1r
VXAuShBmtMRMJ1jHse9hbtgm0XSQd7G8wSTqj9LQ/IdnTfeP4/n2T+PVC7gYxmIIj+w6BeBrShkk
sK9Qbc95sbrvtaEm9/w5wNhbSOL1t/vP5Tgizy2qHbYZMvbtfKkVHGWMgO0qV3ywgefIs13h6y2n
xuzqfrmkO+ub0p3AVKeS4Ppqezi/MJUlDEVb3+nhZr3s2F5zIHnO7QbT4xS20XCdnGJf9Efr5Tuf
LmSe36AViqUSjhB8CFsv14M3ynplaPzJau/BbRf6K0mcxzd6kXc+RsK3dwPeDu5Bes2zla5r+GY7
EizPg6h8ldcenxyG0nCgcYE2AfwwftyVzNNX08C86Snxo86vJu6uKqb7pYg8hv6RS0umYi/KEWcC
07onwvG1D8cs0IyFOKzcvdy/rxAx6yAi76P5+WfGdkKIdvr5eYpLgH7i6B3GTfbd5Q9cd+Pikuq8
cwXQzVabpzJQBOR1/RMtCYAwNProZdb5JYLhqePLRWGURDv1Go46FP6V2tNlyPY2URZSSCuvJheE
h3ncWKsLXW9xziHodqer6RG2gE7Drj+rJneqaaITU3Vew2WuBRHRnJleXsuZrR+Oy7hzkevRF1RQ
zoOZMfzvrxLq/HtRnp67zKOtWW5f9EJ9jYxkmt/6lU9t0fu39l3SUMMEXddFuh+127bAABPJEQL7
FxqMdR6VTwR481CMbITrHmWb9nCl+DDHVLM2jDo3ue9xVeAC2Pa0NTPzDTzTt53MUY5hAD8Lbz1k
49mvpvW/Za4rtgI7ymeClYO+k6aQsyRzNl/WKaMyDGG/Cy7cmJzNti8PKjU0ZhXcHsBwbDFQdnMJ
SGTsLuu6EQZzNGnzof4IsN+0iNFyPcSy1tgppLEM+f+gFlVgcU7wAMNU+WCvr/j2oj8NTC+Y4/TE
uQkKbu6gSFNEQ349rf47XB15kzE/AihBafPgBc1EEUqOLDDreNkZbeiWH8eD5FFhtP10TxywzmE9
lcYUyEiBy4kdnT5EYDHqHg7OlrK754mBd2t6q5YxSBxpU/wleQP3GFwuLNKQTyjirJ7lkH+YBNH6
Yi8HmTAnbgAjOJ3M9xkUrAVznflPxnUXvAo25/0hN2oAjmTwjRLn1LH4QkBZGZaGhI5D0L9aiVqz
S+H/f9TA6mInIg/oSLRuYanumkNQ2KeGaIKGinCB2BEHQgFg8XFRd7AvEQkLwKy8osUdldkKtDZ/
VKwfWNZ1xvFFi1tiAYe+5GuGi/FXoe58k41nlbMJa2tv3rvaGg/coCYz2izibiAe4pYFzYYhCgZ7
r3wDZAhmQVKisAqE2eaAw0c6uba8iJGPaacvbxK2Ifrtt2RYa9AcKBGKl/VXUnWhTLzaze4ik7ZH
gJ38EeEvjwbeUGGuSVomj7QImcIJf6STSmQkieiXXyKLa0bzUMjToeQq5wsi6KMwn6u1nPTdlvvt
c9QzRelBkFYX6950wqcAUkF23MjSSXaSCMXd5dlQZtELMnDcwI675PpuieheVHCYC2b6KD0yczuQ
hAB4HeZt3YiFNnqEMBBWORk1ZzzDsR2LWQP4WT9iWx0vzXrRjnKtim0Paa1r2uAnoZ+IQakqS/t6
19hCod+YFzvaIuc14Y/tbpvN0teaA8roWiijnwskauk1mjd/GIBJHeRsnimsRNRw48INq0v4MVUr
VYalwdhamEAhwcjqJpX6ujUyhmGRi5zulBD7Re3kOEv1bq+9Ks8asx1Fk+HE+1jgT7MO+ss9pyt4
jBKdUCo2B4TA+YK9Pg/VLy9MHRRArjLMOwACwAmKTtBqiIKZdqbQ8pRPk7ikV41TedgIHgTAa3jj
193sjxmF8pyPrI2EJm3WO9/vqXICjZ2gCrNS4fgi32kmb0nVLfbWb7c9X4HfQqXMiEbfxJp2chyq
xQuMuw7J+nsSMqeWttLxmEFG7c3Ey+AfVq8U8bC5SV2mT45h+RRttByjLXEUXNvhXXVxSI2K6HuZ
D/AsWBlukNC/xbqzZDMv05g+DQ1KBbhVMJmLHuAkAlnLHimdZ4P2GY9LFutzYRiyh9bBveR8i4g5
2E8wneehC7wUq7vfqCH4ov5PF62lsL8npVHjD+yKh1Y/9tD5unaYjKyasZiPlkRyTYZYpvk5vg+y
wjsPVAnzmzzmbGOjMiEYs61EkakXVuGd2z7IF45i8qhQryrYCdfeIXStSF6T9uVr1+ialA3APael
G8Nw/x0a7aa+OYBqREEK7obXBOvZavpA4zfKCAdhFxaOKekCnsRctvIi3dlHSrlDPZ17yIPlVKrd
9foPIKqAhAWKlO3Cp8e5I6vDx38va8DI8068P4vZPUHjSJ4n3TTolMiGxTqHnp/lc1/apFJ+k83S
KAWgXosXxJW/es9+uv/a75l9lA72P68M0marC8tlnjDJWks7CVHAoBmfpceB7d4p9eZjPOZMXQTd
Tz1s0aad7uq7lIBKxsQj67veem9bQI3TCMjK+JonKsIkMgE5Ol9/Ndxt5g8Ha7QuDIL2GdLN6d51
oVZheIzdEFVH5ZjSS9yxO0VeKr9esEo+ccVmOZiaBIDl3yjuoXJATbYjOr8XaGEMqrTVDLIxB9pm
jyOujMxkbZZGa5kCExFwDK6Te8gQ3vYHKEgdaypQXBEwMwr69SGbHYYYAH64fJMyTgldSWhty3Ym
0yiiRfvgoldr5YqSYaIno8duOHPAhZe2zxHOjyugepC/kHU9hlc+9VTIbobEVP8zTxCEEYT8yuSa
brXlyrYoIAefJse8LYZWuc7LY5hZdNhv1VPY8VUihTlrJNDYZgNod6Uer7ijUXu6kPh+Msi0tL6I
bJIGK+quJh5xBtgm6eRIP1hEURxjiGkFFX8UaJp2OK0OYsj1t6XN2oJci1AdcU5A1f1Eru/o6wYS
oQN6V+6U+wH8YNa0IO/SYJ+fY0AioeoiXLry2b54p+1DLVJsZ3CXM1UTsjHV4FDSRWbKLO4v8wqv
4RqnXIByRoQhrRZwVt9xw2qzo24v80RDfEN6HMSjrdhU06W8Nrir4rj4EAaa4/6WMEUebYTMrIZB
PZ8/Ub73aHRcV3Io20n06K/zO+sCxdR8O7pp0OsvF3ZcYE7LcDQIJ09XbWbrprfOhQI8W6rYVKMz
5txZQnu281KhcEucxBQagyZB0dn0V2Enk2Pemy11E8fGN3sNqsOpn5gL9EMNtVA091uOCXTuB5Tc
5PsppTO3pxR/i1PfRPXyomle8Ac6uTMDULkVSMcJBNdthYEV9xbgFhrO22pQc1CXWmMZX/zXBKL9
JGRG4yQfbyDusQPWO8bhodvAMtMpVY7FivPUK+RdHKOkHCZCl7TCVDyhJ+DZXIU4smiRuqBybiUl
zgpmArryqc8GDlEIumGcgcrkXcydLREmhgHAEKuBFd108H212RUR59msu6FS88TSH1+pd01mKlsk
iwGpLhN2L0+0rtSUpdwB+y3jJJi84M9Uicv7r1StjvKkJE5MGPq2K67NXrkdljaU5uxj/25o0dIf
iXoSW5620vIUC7HwHUqOGu7n/PJH5I4to5CTiGoc2f9uEGbM1Z+V0OylDtzh6zQ/fVojTigBDBx1
4L4JAEBTjnk4qzopk291iLZlQ0WknTKKX/xwN3nM/hajHKVhFPjDEVRlq8X6IsjVsQXOvmWq971U
8uPsGB7mflx+fR723+0wik35bQfHwvX83Tzq17Z37Vs3AHtZ75ilJBAJg/Um18mYkp2RRe//uaKj
lGjdBZUG00zXW77rTTE+LqFA5x8PVGVYLHQekc9QIASczCO5MCkjscwk4KyVzvwqjjlzZqD7rZlE
F9qmo2htq8MfkQS1kqa0QMxGwLntVrpiEfpjtIrbtQZiEzVr92MbJOLbJR3qIHlkY/EzrfFyHDKL
ce6v2Y3GSjAXhNWDQAl2FkRxjn5Ng45NN7bkm3U/KCahBQ+lFT7bd0qmWPC0rWomThf3X5TcXgnQ
3HK1SG07jrnq7zWGdtIKUCABUGE+Ezz7/lHE5WQ/HK1jQbQ/OS4paq/HEyPAiLn6L8tA3DsvXM6o
fl11HyHhg4nOdZQOJXBCQZlRTTJcF613cZSL7SU4nCmYpx0O/6z/eNLcrz6u1oQItsPhV1DTNXEL
f5TrXXgfJsGc5GLvynFYG9gQoBPMeRmj3Wl8I76K/6cNYpOM2Kdpwy9QBSHAWheY/9fODDvdEcnJ
S4Je3mkuBNJA7dxUeT37PCNnWza+Q5W3WLdcZ//wtfmStL609SWcw7vFsvBJLTpPR3zQ1MDVIxtk
Mkj2P4d7jVrU7eWabdESq8dpJDHDMNZn0GouqsktBqMtD4R6kgjPxPoS0GgO+87osvknj84nRSmn
HCUvzpOGXSQal6oCmXN+MNue6lBTEB7YOuFXx/wf5lFFaD9xZMGxKncRxBoYv1ijGTDW3nL8/ZVI
oyh59rxxDXh6GGhlmIAdXm7oZDtSF6vEJUg7pGEfqS6ZYNjTRijkQ1qWg2qIBedqMt9BXtwfx6OB
Ni98wpSEtaadHt+0NAFHybbZZqNG5WBp1DvJirW9u/3y/Gb3b+9xcK2+4L8OYfyJ3T1OuTVVh7+W
kP9V6E7L6ngUTEB00+X6aiyCORHuKciX6U3kddGq9xDFmybBTgI7jAiThWmJGXKOl0RRI7HwRK6Z
+i5iKd3k1vUK0zGVcMvcrvef8lkprrI6yUTwLr+Cl/EwqfVru/nCA/pGNdd6cNEeHluMzjn7ZISG
0qeIJ5aCQT4PwQ9XD62Ee3PJm+cRLW2Ndlwdq2Zg6azJ5lGyLz/hOJNAeZllscN3eHTGi0PjYgIT
G1Doa3Tfn75PQk3Ag3atLuNaQ2Q0ZODbhCfQVBrW4lkc+6u5b8/8ldR1nRBl0Zp28chPFDPbT1tJ
n31Zey/A2XQrcuiCzIGj1BmZllgeS3FzhF2Ce+OAlQ91VkjakXxnysnQT89pbVqUoFQJsoOubiGX
fU+oXlekP2Oc+w3dwiZWOAxFh7heLnQ+ERFx0ut9N9BcVpCYQjI5rAvjOBC0hffs9UL+sBuapysa
tG2temQSGp21qOYmFcmbQ/jRCSICXKYh1WN5t7geso0q0BK9sPTkMiIJyxg6d4ES9G0iw/n63c7b
ch1hHMVslWRUO6fC9MYGwD+ENE2rsxQ7lxyvWpoY35BJdpkuJQsKrQzFjEOxLohUQgouZPTkQ7Ld
sqRh0hPpXjSc3GiPaWk0UyPHiq3VJU3A7KmrdNw76tgCNRyPGxcGzJlP6X+AzRxvRgEaMPgMohNB
K2iZ4inD+IOvsBP/rgPW+Q8+5GZaqpfFViS2h+igUP6XiKH7ZwHRqCFQhDDKlpOjsAV6bgIgsV8Q
5qIplElX4oeOcCE87OA9w/CmKgoxY4nSF2rqkDy8B+lOoodJIwssF3xOZET/rqw5izRVqCNGZL9o
mfs18txV6MbN4JAyEOaCn9ZqF1PhkngVhcZlBXLwDxqhH8p4RXSY1RKUXBFeJ36eJsoMtx3LhbTM
SPYFn4uwHCEsywVOck80HicJUkyeMeuKY+ZsjyLwLgNpWPkP1ZT8sNxuS/8rw3m7x3i433JE/Xfi
Olbm+Q92iEAURaW4/otXJrO0ZbI3Q79nmSyfHunrUdtw5s21EbNLvw655nv2Q6c4YRdOcRrfsvGC
oa0TQKlUZKJlbUdZvijs4ED01aW9jyeXHnwtKviMJPD1eBKixHhvN2wt/ZdZ6ATn0t18vpQUdwGW
GEjMdloLkFcCH0BY1hrZs7GBBdebC5RUj9FYUxpVfguupnq06Wli3gO7pcT6mqEFNWkYYqHzzfPI
gowtlrXS0681jcAk25hv0M1ukOhMbs5rKtq//7J7jsN9i9dNDuXOxB8cDZUkyyqGXUJrmVJz2uwf
KCp5a/cdbgum3Da29kajge/mzFhxeK1ywl8Zg7aXJHWsDUtgFQ3j7NUJFHq6/dhoZlvrM4kLU8YF
i5NEExQloLhnfoZWv8VitOke7tNj1qBOd8ydmIc3lLZt67QCF633cqxSZIRYE6i5OEvoMMxyUG3n
zAr++6HfusefiHFhIO0npzKmXNRm0p/iyEGWTlHJxnAwgU5g3k05ZxV3aiWN71GgqU+MEeLWLh+g
HHD8JaKX92sEhooluDBZuGZRh9g9s0Mwfot46NU2yzwsaQnvy1MJaLa/bYAq7wuEM5epB0+9hkzU
PVlUQoYnPHtTmGXUV2I9/QcOaplhe85W7V3IH2nunI8s4G/YcNR58uudHzVgZ7t/jFe4tetDa2dF
F7u/jL6o3Cw9YwurZUqQFVyL+swjHxrkbga8+sTc5s3EnHVzX5njAdFhayJkwp9MWgJfUTBIECCp
JrS71ZQRBDflVqW2nQ8gLMiKh6rxwCS/DVaANwZA5p+XtaiGc87Fud6W7bOIgIki9szvIs03+waZ
oCfCz3HvkdD+jvuU1D/f8vRz1/schk4QG+de0XFsrrPc942WhZTqxLu8st4YXlGMu93l8U7QkY/D
qHdWp5xQPrnlbfREHtAAk0aYEio1q9EjlkzZaisuA8p51oMNCQLjAYzbbDDi8/1a/hJkpqrkvhlg
CqC9isdxbStScg7j71ksfKSjUUyoUwj6y/9CYX1k1rYShKV+glfTFCyPQADY9wR8bKNYmbZy80pN
zyxRd/gQ6g0UNyHcSBYWFF5wb8AGkD5z4aogtnO8ervcbq4wYdKimDShgdbHDawlO4VlZjvKZ8eI
lkZJoH2RLLaUnhHWH9d5h2nuyG3G4+75k6oV5MVJ1shfCCRSRdJQfr8kIyEJTJLD11A+2UBiaUeq
H2hpBGQfUSYhABjcbks6MfnStOVX2PMshoZMJCvH1wQUymiG2kjfRFDVYp6nQW7PtdZujs2JICQu
F7Wds3n0oCJ6TIvS+XZtwAr4VZxiY47DCtD3b4Fqh7n5+G8r9KLyVBpuUy/NjAqnLcSb0N6Ychsv
ZOwxkb9fXeuOVbZs3R1UMe55lJre4qzM0hufXkK/XLEKB9Z2HGoizheb7cHktF+U493kl/tpWkY+
7+fBbEmre9+XUFZh0EN3clhcHQsPwBxiLh8qdn0N8vVb+YFaUX/+ZNxKsiMO550sZaP1bix+q6G3
qjheAZzJ1xro7qYLkWzNibHw26DtY4/DvuqfPyGCZ6PYTyQPh59R8BrSv7sOQdYPx4Y/hIQssku0
rDDLi01ECyEWlTt5gYHhWqmP6MQVojbJ0+5QLFxN5LsDk9BV3sgagP9vGzwGhhfxp/h3WqxLi9Km
KRnwaR76nv/ooJe2sezZzTUNPa35Jzo+V1lx7k5CGHKtFfp6NpBLps/0NB4wQq7PyRGcqzS7tp7Q
ZjreHFnraJlVVH0b5THSVm0XpY1UQiA283ZO9nfOBb5oL75HTXekVMbr+WFV7qurnPkPtkkcDzNe
JjjFjeXIoiK1IxKu4as0y5y0JqZv5+1ZhUwGKVYooUxSz4f1bXOs5+TZWETslLXIdr/v9y7YfAcl
PFZdP+aD0gbS0KDvD743tNcs7EA+2rMxH/vm2GgW0Z51bNU/H9vIluYASK8ILk0AnUU6QHPxtwuW
+ZBit62/ZEoVup5gOKQjK/Tu8zkREpmPrT6josG1tE57Do9s3uFprwnxBu51VjyXjz8MFJlWtD70
jT+wX9SCSJcQlLOrsEpm/mfnNeGrckIm5d6o9zVfqd+BQkoSdAq6Jf8FwFPOwDYFdQRvY0ienRc+
JMwg4dye3qmxAeGkPLa2RjZn46DbcFC3wT05cPMQAoduA/xX28Kk4OpHHD9c8Q/PXd/8hccNdCJu
sX9XCg+bTTGYg+/hGxPvsS7OzfiTiLXoDQ52ss8tydkFakf21MDtEpV2XbrCiLDDZP1opvr0lqtE
JynZL5aLdhtuV+jx/h9HW6r9tPmih6H4KpzI8Zva7TVWkRS8yuWdYfjS/0iaT28fmx5QHEQ1pPht
CeO3XVFtgXmzbYQX4Z/znUbxnfblwP7D4EBquGc5BB/vbNLmL7w+XOasw/579kAue2CIiKmqVfky
4rXyVZjdUbn9PA2pCO00S5CLMM9m6TZD+P9kpO8/icBjoByZJ16P6VrP/PcY1f+SF2NaKYTE2e4W
O7t/eKVzRjgOzXNbDVKCJXzo28x0IZVMRHurJKLnZIMsstgHkfHO28m4ulWvwnvibp1hhl7N6X3x
VRS3paHA0lTjMRwbmy9QgflPW8K906cvgdazG7h5T94IiTzSmv6DMSdg8joHsO8zEZLXhzeaYIbZ
WLg3YJj7NPZWWpDuUSIH+fpBqPc9KfV/m4BoCFLB/Dq5HZ18HMa0WxdfdWuR+Qr8w8OLvoY0yw6c
mDmNrUeQfGbrGIjQH7tlWLkTZGj5F/gtffW5W2+W1agoe1kTr+w+/yWjjuNp4cjIxKnzE/TK7YG1
brIhVlxpvfQNX2xWzmSLYTRc2hnFuE5jPhJu/xBxEVGVniYcfgwwm64+xksC4kTpA8TFSnQ5WNo+
kThfwfh7NmjorciJ+O++jTEZIbs9T7NDwC5lh7pyQmNRwByKSi7kwdEqQmNfZw8VTvSOPkLiIrTU
ydKYBaXS+fpjFmylsYOQRgJzhzulJtMWjZ/HDvvTFstqKnAl/VPYy7M771ODhMtlnFfFEnvp26j9
NfdqLemcetjYE/kWe5TobpzFFk1iCD0onc//M7mpozF9CMxwRzFsw4FPlg+BduPkRPxmIa31GZFb
5gXJz1KLVKW3/vF/oB91sSSMui4RJo11D08+D1x5XCvRvQER8uzTURYia5LS3VFisgZ8CaYnycvE
ZlgEXlEK1QiXOazjvXCa+18lTkHTFnPq7AQkhO7iUhEhyd2LUZWPSWekxFuWRUmlL31ZAr3EyejZ
aMW4MmiWoHOxhblOL1RcOzwiKF0Uy+UZ16skWWq3/BDdHLff8NpZKDzeTzp56/6An2UwwDbjkb0F
206Ib2nPoAgmcK0kd1QJfyQMESObu8yz50+Ip3/JDsDJDP2LUK3QwvqRA5MqOqlnpKm8ML/ggXAe
EGJ1Vd/8/9FlmrZpYc4fwoQ6toKyHx7GStjfW291wHAt0KQNYeiDTXHY3DI5m7QTtnFAni6XeJeO
0WNiii5I5MShWRXSS/1Q2KnHnB5F3Ic6AbJOB2Q6gM1VD5uhr4ZkFHX3G2xDYGT3XH9+pAbnc1Qu
MUgxPtRA300faEh32Ay2BYY+f3EHNMVQg5dbtH5211+MmOgaTfhGDG5+NbayMuBro+h8cbvD1GGN
zhn/TB9ff+IWV8xeHp2GMUQCae7LcpP+wrE1NkXkYycpwZ4uJ20nDiKlml5IBgdLB9lcDr2FCHmb
k3WckDpK43SCwldkL2f5G4+zsTbxKhIcsr/GDly7s5tlxCsSf5ylFPk82JUICM7bPK3SNNW06GXA
KtS6E/bsa3fSLG5v6W5wDISk52rVN6X8jf/0dHIZOUmcTQNzPLLR6Esl/RWSP5D2Kp7kKl9zOZzz
p52JcpLrrIRhohro2lUrEhVQgRx0OOzGAOR3x/zTv8Wv+P8XCKy0H+/BYdbtI2uOMLOryqQasURb
xwYCrjkir+OAagq/If+TtD7GaZ3naV+3JzuF95FPlMrM2GBLAg/Shwdlgh3SlbCaUVIFwWpOpU+y
2lnYshhUL5yIPenHZVe4nvWe1hvtjCKY6r7nipSLSW8WfA5eXiqfxffrtR2KW16YP30BMBRuvYwp
7pTrkYn7g/bVJ1PVO7DeUI149uuUWm8fqCQG/FQ4WuRKazO6ENY5Wd+rLIa93pbZutxpNQwsUe3f
gsktZ+Gs1m3mhv4DN/yCYO2eHUPu9tsK1z7l+N4yPGFxTqIlvZIjLQQEbZF1wqAvAfhRn+u89D4Z
zKSQ9BBqWDm/WNYvhmCzwLvb97p2eQ6eFVHQDf7Wog4wuaCKlRN+qiuAzNpqsDGHsdwVFPitWJI1
OEybNEHYzv3mkjpYWI05ydVAWzVAW+SUCbu5/QHdmslrV1EikQPgug2ClkSUAxjeLeEfbFcRwvlS
5MB4QbvDfCI/FV7FS+ilbX8pvPuwSXbphEDj/atqxEdsPwVvsNVHWG5R1wpD88csH89g3YzhZDkO
IIYvjjwJshOt512hWMp6u4pE0vXdpD4HL8BmZ6IqtOKCFpHjr4nEL6w4/wADQtBFd0AVd3dYD2Hi
hpMM/fA7lGWyDApQZuO/M8VtnUqNVf/EIWrodiYnwyxBrqdA6RaG17tp9KMhH2s/DJmSo+jAD0Zx
7V3lV0MC3nMnX8Vxl+yqetgAJeXM1CF2n/ghp+4Yt8afiOfSot2083NHhKLdJFmO+pPLRXGViFzS
SJHNuDIbfhcJvigjTzN5DxZhGyLE1Az7p6j34NO81bEFLjjVxUqGwjXybkgRKKtkwaaPAgQRmMuR
i/Yk3UoDshNpUIXUmic2vrYya7IBzAgoWd1kdeNk5ct2YiidQRDOmO14lP8ybK0RbSxfveFXXa0x
qayXNohO7RPrmg/OcfNrAWO08d9vENP6rFGvbernc1LGUgMpur6hG/UQtZ7dD4DoAoJhiK2tiTyg
CsyMsSba6eXFPXOzGq1B7ICjyu+QsBByipFWztKiCjWJRYZUaiaQ84i+aNMB8fT1wuFR/903zrBX
8MB3Cxpy44Ce+pJP5gvJspvpMlQCI/aDKfu4tpZfrVft6dA8GHQeau/mHwVO6OE/BW1+3xCKvH0f
Hvp0l6odjLAQgE+erbBvN85yFsrUHPWcfseZksOyxqhk6W/VJIjc67lvbMYzgZC+FOy6YAxu6hP3
Q61uz3F+ohrOAUK/yzDi/TfonqEIIpzTlnFWSYFU2PyNH+MbPtE4hUwurNMQepJB7uGUPwNhT7fy
6+aWVylJnKQNyBSlISSPQ1GvOxPc/ZUN+N3vQFx4u+DwyAgaMJsTw7ce87ecuFI+x03Z9QtB4KWe
WESjNYwHvRpNX3zVMFPdPBro4nxxP3A8mfzSmWt/Ki1pTD23mAEPi5//Xw7Am6g/4NhCSUN01e8G
5sKUiEHwTrHZOiu3Ok0k5fadTySQ8LzcpCp4cuBsh/BVsWsLfM4EXK5kBJk8I9S1Ctjeyl+HH7MQ
a8BB8nCjI0PmjgC8kZHGT/9KkLp6dbU/jL6ZFMSXLF3agpY2rYUNi7sMqZINKYq0goHdZyRZ5Tjg
YZ3XmlplX8hPn7bYyPp3HuTHt0/u+9lBfmbiOpSrh/5D/lF0kJANTyAeQhEA9s6OJNWIMfmN0A4a
LoQmD+28u/BaC7KLa9nC1qroHVFlnmshZ7kYI5ZnxLRRzgAU3+YT2l/n3A6BRFt3haD20U2ez1L/
lc0MbTjwKb9F2x3Fj9swLPsuRsDE+cXLnmXGFsqoCSeGqhI3J/M56sS4ghZu9XbOsPGHpyYte/cP
qxLMXYvxuaFYBPuwnVkGvApff5w8X+shR3gqshViZVklC8edo3gHJ2WxjTJ5EgPTwG0JKokVCYfh
p+eVlPhR3GjGsMipBa4Bpax8Mb8nY2kKHZSssFXwn0NFjJtnBqxok1G043crVD8xAwWP3M16OsTF
L21heL+kzzI26NMTQsX7WCUvbt02RHGk35SMYqx3Ju9pRzScc517YgW/xradhmHdPhwGTkaQIuMY
24bZniLQNogJKQROGoMX4N2rVVe31EHUgpG+wlIHSX/KDlcLB2apfxaPswUonw3WKpS8vD6dAiJ5
vCzgP/S3jirvPK3FpLn0Lmlt15O3uO/edwMDCrfbzKMFRxqFp5UHXyKWVrLezrIKkY5INhzuEC/b
RLbXG8vC94AGe10T/sVZn+Q6QVFkGp1HgB3K+oMb0sghn2UulAikM66/KzwLeFfXPnwvdDcAj/w/
ENn+WFmTbUzL9BtYqSVMKhMOsghjdZO5S+avd6rG381SCNcpCJ92mo6SRFB1ff0kPmd0zA9yaWuG
zShlp6OO1wgZQ1+T8E7qZG1V6gw4525HBmOK3pY0YAtIcyQjQ8BnUmf0NW6bihmSv7NVQfmCWdw0
7pahDfeWuUxsdocgd6AwBnFQWKN6VFKCvGd/iupX/kD/Zvmx+R8rf0oFDX2bGYBAAk4KZGul8tWq
xkLuocDONxmjRvzr0JWtC8gWJil113SS7An5sZ9RX4kYNUq9RQtILrzrK+TPnFnN4z6194GYLPc/
4EjvXaQQbBxPTDWN7L1B2iwMbCR83Pw5qYzK96SnfgMALuHKrm8fXDZvFx0+OFn9TXNPzyl6TPG5
dM95iwgVPpUGEnbs/408ICGxHknjWQ8aZkMxfq1mBHR6xJaUYAYQhlSwq888FudNrdOrGZuy8IsW
n5J3HEj7dcWD5SRJIXmBh2XGMr4mRhcgC0hJEkLzKPulRqkVOoewod6WknCR80O+cZaMirhEtMVa
66xfUrGT/m4e7igaWAHQZoJVIDHmZ6NFWsD3VH5gNyB3CamgjLita5uGaUgfqC3SAfIcprGQ1io9
IvDqnPmwWslC0bIqB3C4rCIooddw6k5zf2+DK5IxFsjvNc70k4G3R9s1tsws3yjuyfHHFCpomPqT
iewsPfD39g+NtkxV6q8Ii3gYU7aPJBg3eMTCxiMCKj70pxEHFXwtejc6cUVUtzfGpP6nA93Pz9n/
E2wPby72SVjZD83knRwVe1DfJp5zoth8NRoyLgEwCGVCe0z01dW1L7LSrkec5uXSlm3KYDu10eA6
yH/a5ID6aeAEUv9taSPku24tRUIOL41zbkkGJ7jYuQEddlwwEZYYoUP9/owFDg360eZQlaS9VSCH
Zs710z0SeIbRCtnchgV8w93Q8ayHnfleN0Oj1zKyNkSjHQ0TqXLPrtNuqoiCvEeHJZbZh+6J6gA4
vwyk4V9tG+FG6prLUCdZkgi/P/t722mpEEliTyMSXI1gTA/Q6mTCNtuwcGwTKiG5pYtQCBVnQEcF
MUs0rWhjwsX+NAP08pRIQqk5yv1amtvbGIuhRAnKHj84Csuf86PqGiLW+laV8DEzSWvgxCBb05lJ
18Bc4iDyumOJzjxEY4x6aehf8SAkFAY8ntKOEbXYkkkjZTUHbQwfPsEw8mXODhtbp04e4Rj3lyvS
swt5ex1WP1CtAhvMWfflFbHbFDbhV79viAEQ6RfPPohxKIqYx9rSKltI6sNzuvL1n0irqxEGSalE
Z+YA0IhwXyX/3Ed62fm1JRi8+IG4A9/VSK0GINO//SNXnrN1rJpxkq0R8vNzFRjpNnKXoeiM5DVi
4I5oERccHNIzmAnbtDGX+XhWMXzTi0EcMQ6u+/FUNI5SIt8Lx/aM+TSf+pSzV0nB0NC2oQ/30Fb8
Cz8a/7SK8Gy3rw23LtXrwcba1bPDfbeX0z2iWEV9VwS9Eimz08l5epb7Td6+Kmud2VqoFckYFSNE
+r7CFEZlbISgUvirpy9VF2LpFhg57AAJN6W9g4hofPIEpB03HplFMOFR4aXk5p82u8wmKWqHqj6j
kBZhza1X1r13nMOximnx1aRCPtzfWVA/8qVnol7uDyf/oNiK1NyYPPqXqPm3RyNGtBZX9Y8NGMUL
rCl+cx4OUsoh76DqvPhgP85MzMbkMci0Vufw5QGTmy6d9Z8GO9sU4IW4WRXNxJIDz6Z9bgczUgRl
/aLW4ZXwlPs7MbxvYCXBh/Oc+qvd/EemJhhviZPDn4zp0TSrcGjlSzXiAn7yrVCyTi4mDRaUqI5o
/TbNn16oE/vMM5HQ5ZflLVsFmvVoKY/owd2uoUGupyZG2bZPrVfk6/L6Pgd263qSMUH8N7iEHHIh
Uo6hqJ2BX+exgBkDEOXt6yF44ZMC1pDmjjUpDv6Nk6FhfXCCEiHwJPIWNy/EgiTu7soMGpSyza3v
OuLKDLK5x0lfKdU7+Q/+RklDCjF7O60Urk6/YRPJee1uZPfvczQaOoLue1S1H3NjCvbGZe0zbZ45
2oOCXyyabKGiVNK699s3+G4FWDsd274byXte/JVWGfTJo4LZ6G/z5/4yBm8/ODk9q3rOG79htbCg
etfkJ53v87lIFRm6m1dcbbSccj92clWxmXs4Uz8rQip9WVU/WT1QwGoXw00q9uYbzR5gs1S3lSB8
FORQxo1fKK3pTkf0hW2adfetVB25xraOyq1dVLCOZuYn0mYRrZq5F5Wn+9v00pCFzglNID9Rn0Cm
2xqw0vY561E9gYO8CxUgyWOSvv2AmmGJj7jEyNVEJEigdOcoI03f/T78LmmlqMAphZnwXrfa2W99
NScn33umgfG2gw+9GzBtLAzGwoveqkKICBQq6+I9w2WHm4zjdHS6Tw/r8sa72ELjD4o3XUjqLe+T
hKxLqm+hqblcp5xSKK9jhWaz3B6Iz/wU+FmAhSYZk3J6Ey79N2iNLJ5zvdK2lQRkUrzI2h94xhbf
OUOo/zByvUSEo483QrC18/APo64BTuBQd294O5qAX5KOClA/rS/D/mI4fLejvJ8GmtnzBiu/XV9i
0XKzuRb2DS7JrNBr1JUk4xpQ7jCMqQl+DXfzejzcyvZ9L2cuu22ahERkicrpjxjJXcU8lfcQmNW1
WHkcq9Y2pMHF9RmOdOZUm2oqaB7hTobFHWJvxHw9QqS4VDeDJ4SDLEmGMGQVp2XqRkKz6C7YDDAv
aMjT3ZB/11sQP1jLsVcVjI9U8CSMT2uSuCF9kTXuZXRHJnVTREXEy9E/AjhNt9NVACoCZxm08ENB
pD+8kX8gQ42eswAbY5HRNFiIdaDkX0cpDFDjXICkM2dktdp0RSzuo2npgYogV4AQ5jTvq6sh6n/J
+nGPnBMj+sbLWY4V7yyv8i5BlzS1FvnEPBfPfWPD0CWaHTR2IFaRR3b+8EutqCqTlmqjX3xOy5yu
zKoxJSnkoF4vl3iECFj1NP5jjMmUjDoSjr2Nao8UJDRW++puxUq6Fn2WdbJIVIBSzf7XXiRblMH8
PgB7zjbAKxiwSrtTWwzyaYHK4oI3P/FXJlQ9yFJYWhnYG+f7pE1dMP89qwO6CRsLJEmBSiYVDIWx
GyDp4gAIAoT25H0vhNs/J3hC0IeEpS8TMw0ias4wk2UDOVYU7NFWdgGtHObB//BtdJkonjYdPbQS
YzIVfLgGYEB1+4xdgET2cxvtIGD2sBMc2/cS/5+iZguG8CohujYoYIDarodqhM6bmZaM1cQzFXqO
31j/BkXb9Ypuv8kvRSuoxVyMmGwgy6q+osuCH9UQMnCWdjiDwRTFWFyniM8/ldvN7jiT3ZNjggbY
/toh2rkS23FO5Dp8s602E6NjPYXgHbbVum7VSBu1UzrkigEVNB0EV1VnZVtOCgtby682Ipww/QkW
x6rUTSwJ/ZC293sE/Ng0sprRWyN6TVHvd4ztPTE5tfMnUi5Oieob/hgyw/gylGBNDrRYZxCHHs4S
Y/jMsb/4pTCTct/6U4XpHweSSigy5ezUBhZCjffxroJIJouMkCgmEYEqzToVMgt8OZH8aGmpJA+l
LsO94qcknHJpj30byZl59DahVCVVKO7zDOxtN1ySIKz6PhPmemcBnMncUyHCEtDhYhqpfQkcD2iR
9qXZvnPghwq8/poAzE0tCIYa5h8kM8EaLbV+fhZjqZTuhe2+hRe5RyhcoaaMvIEEr+N0KVhv8aYj
LWvG2CJUVizTSFy1CbYazkWYUQVLsCwArpSh9q0yZLd38x0vvOZRPZhTnpMzWILXLupQppBwV56h
yh7S+g7Z6V6CXk6VFREXufJiuaD21sAwlyaTDWZ3wMmJaFDh4LlNwCAIFlunPTPi4kfAP6P/3BEY
GK7i2h7j0mMQFzIIJARYZdQ6bsEC4i0K9zoA8ycVMNgJalADDZoKKny+AbzYlkW3WZrGGAYM9LNc
XYr27lC+Hcons3xNZKZswtr7368T58Z8AsogQTLSfmM1W0O8Yfefqrww5JT3Vme+Av+iyXk4mMhp
iQtnPEEmnOcRqAZ/qc+09I3kua9pouWtqyNia60X8GaKhmEq2txT4gCCfWo5/rH1/cbDem0yhY9A
1OzUAhZCeRHPmOIgppaExFXwpJ9MVS4JiAD+Lu/0Gr8t+OL3GMJv3nf/UWKnusZXqZTwBlG2OMAk
z7EAbdmuGB06f7yxsZv/BOxvG4r1ZcvuN7IYiezPC8wd52cSSnUzaYT5zT4iZUll44ifDWTNT5XE
f6iQ9BCyk8p6MAdXZ8uSX20ko9XRXE1wmhDxKfieqyobcPGxvqYmcKIrV/MoQecYz68oXaFsBepG
d1tn6d+wwGWouqMxHFxb0STR+3wkQSS/NGg8RXj3fe01YIF9FvMctBawIdp1v8ggMXKZwZgcJb4j
KiR1nRCUb2vs3Js73FWMxpf9kxn4vsllXQtFuIkWwyQ4yYHIGW6iArFmucI/Ru4dAADVOOms+5GL
LHAguiMqS9WQ+M72eTTaxNC535eTGwFE2zsl407JmelrFMiLCOW/c3VhEpu0HNg4hTeYTYPqHymQ
K5a0vDkE4JLYacajZMEKNDzIW34yhsxRBUrJtNiuHmlW7UplyhKOBrUrkSmpmw349WON8F4xV77F
6hTHAigaE/04Iy5lJcGCkhtFi7eQ79ZybREZOYjr+Ss3Vc/GuG2Fvj6k/V3xJ2Nupc+q3/AVl/hK
nN4Lwn+BW1OiZTN53of7uSgTp1x7LDNvscaT/GMdTG0Jhv0fjcWr70GtcUPnIwrmPkFjUSilrs0w
yFatgRPddCaJRqzh08GZ1ezL/QB7cnYYJHJSa0xlCK+//C9kOtXcKKXSuexewT6rrtei0qDH99GG
WrWEjUMOCr8d97pHEv3iqiGroOOT6SOVPG99iRrURPUa1+OJ3kDPPGj8NDypRnudsNPBnAtGTWuu
37L/Sr7hoJ0dvd24hjMMTw5s8TR0n8AKDBv+7gvD9IN99k8OGnTBVrRsKTBJX5+ZBY3UDZoteGWM
86VJ0wXaDbjCvNp+CpYUpJAR870dSRToFa1cWb1l62sW8XyKi/hrRfQLohkaAiJFDuuTDPyRPdrn
SV+0SWTNoHVDSAtXyiSFnSnkgsRa6xhecwDofEhD8BBxrz1j+qeg2s+IbsYP1cEncmZ/MIMBuemi
B6srYO3sXKOQFGcnCF+WPf282q6GsSPXpVemENz1gghIRrbW39VkZYDMm7/aHe4A6+shwhG0DcVM
QSlgUjCVUYF6D1FDyRgQns1ipHqvSJgNQqU/1t8mnaN+Q68uGjjA5c8FRto5++pycZI0Ux++t8Ch
vujgaMCtMdR4US71rpbzLtwy409I0nIBgztDINMtlbb+FYnIhT48cw+SPe16FkZZnEUeHkbqsDZ+
5wruCMgJOVTCMm7sk5F+5laIjtFCWqCQqeVpqG4HH1PFkPZp9wlcbc376y7es/Dy/yFeO+Fe9UdW
JnXRf3zwnsH6ucbvvx5EyQt/SbvpnJ4Wrxt4CGjGAN5xb1uG2rSia8guGsPDcLkZhIpTtcAYM0fq
SwmFmyXWuLV0mMKNijuTE+MWlfxRD1uvdnKJpeXZf1eh2y2k0niA5MxsK8d0/jdcZgqBz/hX4hlf
U2/jyYjhJi6pv7FmLKTnHQpNI93uELYPvUt4rQPf4N4PjX4EIQEizVUJlDhc3npQZXrfE8RLWwXS
xa1PqCEmdcr2HAoLYoWDzICpErwGJ52BCPSCwZgaytM/e3PC9qpyL4XzXVjK0D/4Lm8ER4WBoKLP
qZvKNDORALTM1Q1sphrM18dSAeQw7jnodKAi0NzICFyufwgLefJ9tqaMy88ZBHxnvAj97vZHm8tL
XMf+gtxTV3uxtNWjiIU/6pVItNdqsC99FyQMyKB0n/AuK/3xt62pN66kxO5sjBzQz6MrBmaeN55Z
FKyE4S9I3L2X0eBGbTWUvIyvGhNiEz4N/yfuByr2tJmz7+1nBJvHRPhBMV7NKgmDvZ8A+dwum7IO
PrsTLkYdF7KhZUycKdFtN7jpxeAhEd/iCNBCeVyxhgFdF8mME9Kq9uTRi23mOXj9CNfBAClDbMSY
+/cHDUivwYllK/xvHTlXPZ+sYxDMRsQwrkG1YXoi7gNB5FwAjhKaXo9rc/Bl3vNsXTHqkHmZyNHz
a6P0MG2gWUQSZcyrU3GYp7TW7rbomYUBVmavVSUkzWInoKgZaF472dAC/BpxhMaSO6ksqBQDfyw/
vphy0CbD+Vpv6p9WTuQtfYtKenqucAX+OSSaFPW37osIKWMBCrGNmSiUoxySjNx5UtjMlG25qTtc
egYCY8Whj6LsLcSn/IipxzpyEkx6TB2/ygr6k/ifwnKVtbFbtSypZc3LRID+YtufFt5frfDHd/Tg
ofgT/R5TL25SDzW3WSZ/BAfNl6oxEDlLVH9obVlNiM2OKmTudDyh4ZJ6vg96L42IxCK7MMoI4FAX
CRjbXaAePdAVPhwAEKUTLh32TBEJ7+cGbzXMjplEGe34K1ujXqcHqKaLjiztOy26RV/UYgQhtugF
PHwweL0BwcUQ2d0ql7YNDMX8vY+0/uGpKPabBthqpWm3wCZCqRFqT+WAwTrtdtrzjpG0CD7rGnLh
p0SbGcHpaoRHweGzuyQy/8Y4rVvs4wcTSeWjVNzfyfRmfVxZiNr2WutSryVj89Zi/uzYYDWeVWPb
5xablLNKr1FztBDWYCDGytTkkL3qrqRYm5VWSQ+5/omQLVKuq5yvjUZq6N3NYlkziN+1nG2hMPbK
k6dJ+5y2ctuAIvdL3p3X/u4rk6842UAtPvR6hJGmM9jYR8MLFHxEU/rrG3HbL4O8Cp1ZhxIgIxh9
ywfeFFPJug4DeDLbi7adK/0k1BdBzocrb8escxNFYOxs6fHK+iA2jj9NY/5mtl2fnEYK5W+vx8H0
CXEPkzAaQt8JZoh9QqEn3tdzE8sGNhltTVCWvRIRAx2EFHWOkt8dvJhA+UL0b6d0JiGGefvvKdxx
2wlyoK5apgreRy5TXpYKTW/P/wdy1sVNHQAg0KhEhY2hzb5MMLwxrE0cB0HH9soVg/n5dwsH13H9
32LNVhRy4v3VeL3Mdw6qbUL5A+s3psFt2kIDDH3/xbrGOevy/T1C960RqJcv9dD5/+ZuB7HeF45J
l3cC0p6ryk1s2R2tCmRIxy8Ftab0pk+5iZTj9t+hCyvqEGk+kJy+FTTtgr26eHzM9nL8f9fRDM5b
S5096SqxHuFnlcIfIWhFzuKcdZCUgT3Q8gHoG4HDfcEI+TlVcrQC4EZoZjW5IlY3vgem7TCP9KI0
hLy3nnQ3cOLKKgvIzdnTwXuaAQ8HFSd47SIy3Vz97DwMDq8rIGRY5HQSoigQ7Vt6CDB2Xxly0my7
tHJVO/F7+QZj5uupFVwcYike/a1boveIokpofwl4GnAW673Xm9Aha6f4D7O3sbGCqS5WP1HLn5sK
mwhtyrTgS/FzpXn+n0SHdOe4yEaChsaZ+1K3e3GW39FTYqXfPvkAlEIAQ6TWEQKsb70TTHfF9kTr
QiadSgiQ32Oc85Lp+udKcodP9RFef1Dq/S6AJqlNxfNwScn0cQpl27pHGPPNYvsM8vR8oXliCPYH
mDehZ3ah2wRbBiG7+R2r90gD8p+Dds6wtn79W61IZ8p4HWDLVKbLk8rfh3c47Ytw2yWVqEnkjJp6
Bhak6Y2K0M82pZc6vfILZ5NdlNYEynVcETd661J2jQBNs1fPH6c4GvLOtNsDS+HL70kgdwc9iCqw
kD/z88fVIweWguZLwpMSD3dU9dFPwG9Vrib23I4inzHpgNrvF2zNq5JzvMxRFs1YuZn6yJ60KsDj
F3tTt6GkAoLOzKvwLgcYi2819gGjBlzffFYK4iwT9JWnq7ZqFXUlJjh/xSeyyPIc2Qc2Q2Q8bTUU
MbrR5XjIvZ8OLzCrlHsT/iILvKkZt33YpdHGeJmiWE41l0qW/kLpdN+x5wZ33MNGVPwFk71VNvd4
6G9j7YGMQsYFDpwIlr+Ep9DcdFmVY2ryH8McQKfe+nXtkNDqxtfL1EHvFpPBnPt2Sc/u8SA7nuJk
C2pFwcWsx8g4ElyMU2Ul3k78wMrnX59z6pc50e4uoUn5b1KSuCdQqalsdmGChCccIQVJVy2Nm+9/
OtBWZMxtp+nEbCtReO6CBZfIHdoxWRoCkGTgrK3neg9LE9AMI2NY3MJZFA+gljS6hO5f0iwCP/XK
hVIBq3OXJbfzEjVpd2W5H3L99qvugdfO2UNMGItWeLB+a8O3ySQqAuxjvZW2LElxTDoWBC6AqVNs
i0E/wlAkk+BbZmah2LzM1WnGkGlj3vmblX6o2W5ODxtiGpGttJZumpoj7WdUw11JCYGOic7Xen7G
ZMB/FBnWGjWDVKL7iPV90jZtZT35/L4+a8/tZI57KZwLpqaYXfkHFDG8dTkt7QbfqUPcAg/b84uS
7WO1nDsLIgvFj5nDhjCpTQv4puz3CuwlJbonyrkHzIrC/FVzwdG/0a2G79ESiVQGON0widfbUosO
XtBZ0IY8z7sv/rAAwdOCNkoEoxt9Eykb5WuiIACH+TV7xEbUmzoMZlo8IJrHzplf1noVvrFU6uA2
7sQ3V+nRA8JQw+xcW1cJiv0ACY/nJ3fdxxV7fIcgecS4YT3QBjAPfmeGDesIM1wuiS6nTdYwTkrt
7010ivZ+jmtTTzsqbCaDqetG8C8dMvX5cH2n0rCmDvVg9ykTn9SVaJlgvwtEJZ+iy2uKD9lca8Ca
OdyGMPeWZe01dsFPm0nZ6Wf7nHpORdpM/dXDVmgK0VNW6AvaAgH7U0AO/S/q9vDKU2JrKHXtWfPo
BkC086s3HflugifqilyPk/f4Uz1b5Hj1p+jHz35S41dS+8Dd18FmEAsz3cyl21hlY/1+cbVKdi5f
4QlH63Wf+E7g8g6I7yqbasTCHBcc/fIKRUlNC6DdjuQ+go7LqfE4Ugf1Kk5HiiWm9KCP0NVOxQ5E
QOuzAlj5nz24THS7gX9sR/0wFy7dKyRxc6HMwoTDhef0Oi4nf+o+Z72FvEL7+/04qYVCjLNT6by3
TlNIImXCLOrmCckuog16nzgoch++XOfxlOgMAwHUdJ6HbSX+4Z5GywerNwQJulwy/vaUuoW6QXcm
8h/Casp5+YdG/syFMOKko3/N1kQGCARP52DcDJGVJhJWnQBFl7mQ241P6hrWAVceeFw4q14thi8Z
HE5P2Q3+6wBMkNlW6t2ppsUk5970w4Yr5MbIkdghvPJbulamXeMg9AQhuA7sZ/p+7+qLbpqG6yoI
KmNywkizNY1fahGO0YOMdEnN8ItiU7i4D4JWSBHjKT+ZuHVyPPKjoi4BGxcUhkVMKK9WErvnwizZ
YH/PzDrw1XvcAZQprbb0Ecu5jhH74UIimO+XKzS1TgsAb1h0q0qeSX0T2HJyTrhcNIaLSS/jycwd
BiFw0AjcFQr4BNHsWQThUaCLhz1D/aoPxbwjOB/8UvoR4TiH8SH9Pw1G8Ki9raRbjH4UhlzcakfC
RsmcQqqgRxIpp0Nnze9XkydHrODT2M8OiGFCVgaw6HKP42dI7UNMFRs8e4pSx2KyU6nJx+kNy/Mp
qu4xsF8Rv/oaKvjbsX8F2IJwS9eXiYL7Z/U++YjmelG9gWuActFmhgwKJ78+ZtBwqNkoJDq4UrxM
/IxpYDT/Ju9ApFOSBPkp7lET2SkWuI+SCN5l4dO+p8YXSXaXY95Ysg35pzUFy9wiA2U1SZ+YpzEA
CL7TqrqnXyw7OFcqQjMjfkrNsKXv/qFEqZHNxt69vjyicf8106S1F2XhRDAD7zxEK6jLkSUYMQ5q
ms56oPdmzeys8JBddjUqk5myCXAB1bE901mrjjALa6NDaXhBHIIoBNqWNjUsQKeB47EPPWwUE3GV
CGowoZVDdX65K7J+rEiuseiZq0UD6E8bgbapoOlXFYB00QDrsi7U63E2wkmJQ/U+rjwUU5GffJ+4
lIlq+tcPwOeeW31XEfPkHiU16VxWk/Vh6KHsznUwY0MA5X9iTfV6vUWoCYOWAy5niFfHkD3eOV1a
sAGLgqjswCvi/J9DNDRI5KS3TWUzZfXv8mzA4v4H8J7IN7KZUiagtAVJh2VxCQjj/FMf5dG87/qd
QyQts9LuJF1rOOVuDksFp9VXBstqtm5OAo/7QJwbxBQYncNFFiGZLdcAPlgdfee/pg7ktUBmRvdq
KWmJv6CbhtgiSVtEquYLdveMxhFUKpQQqGTgPmSBH020/cdvxvwGiJvzYavRbZQPLwzvxJysbSil
MDkmyuUG4T/8pyCwM305CUcKQVl54YbToa3UrYUs8fhZC5l6AjaWnqNBMslY9h8VwOQMhV/hLItK
mGQJiC2p5rI/VRRw/vObTC7ZLuI8l6vkkQ+M+9VCN5hJ2VQCdN4d+CODBuqgB+7bG7G0WkJZOIir
AY6W4YNAlOEOINvKcOkCA1cMvESwfN/vPbfcMqHWD0wjghxHMMZ4d43oLROLdn8sSq2+pkAmlVZK
W1qkBzNx9xCn5zTutvjbNFaNZs16opu0qt/0ElYTZILNuL1ExRSuX9/GlKuL5rOaD8Sdcm16GhKj
G9p9oPmRWPw2C9pahljc9nhuqHOrPHsx1ucaW0CNQyzjgW+0ekGYrFKrfRtDRK9r8boE2IblbaDV
7dK/rzrBjT806zincmtGKlZX0o0yooCAxrKZgUvIj/4Xfq7zGzM9eby1yvHt/QQy2coZTynQ+Fth
2u8BNAqq/bs7YzjcsECHblEel90WtYk23XBX+YesiKYBNe+kCc792evmOPMu7mKvLGig55RZqvBN
TVoIxCcK/LHXqEwIXo6iKS41V5iKXhJDDKDvKv8rDmDQkFBx7Rs8eL7YO4knpmHPZ5MtTXqjM8zs
0k/q2d1kutlbqz2r7w8YZIpYFRs5wcrfJr69cjx4VHZ0RbIpB8BqFgJqmkph0/49hYfUnJIsvjcu
cSR+V+6SchN8RWwf+as1wLM3DXBMpF2zSmbeSIaiur9HIiPSQpJnLwjPUV7G62Lrosih+Q9fElKT
9loIXuLqsAGVick+y6djZny153pgZsvjAwved+SCpWOKaXiZBPktzuDt/YCEtcDoSxI3xyQvqKas
suvk/00ga4LQiK6UqgiUH3I0SQAIeNkdRJZUtx5ItlFMRyvjsYha66ACXt6Vskgr7FVtzz8azhoB
1yqJEXpvjgG7LpQgm9YjYmVOQByWx5nuT1683ISQJYyrCl4B5XM6IhYppUBngF/051gvSXWqqtsi
dRb6CApBKMBJ60tdaxvCOXnwpilS/5H3wkEG7d8NSRyDO85GBkfbToZh/+OcCX4bmlVFJ3rxi53U
5T5nYv2VCXol49qn0Tc7SUdrnRQ+uLwAmHJfKaLllbrA2bsvkumhMFpWl/lE2+r++agEs20nj3z3
ZLBR/f0KtVokxWONQSqJV9ZLBbugvlYxpqp5SJNoRUtdkC5xA5P3gxiApZ+r14fuSsIVOOOt8Zsi
lElt6K8YC7CLBh890AP+BRWpCRXvitPx3CxVTjb4BSlsPk9CwA7ayJYut1BukdNCuwuEM0BlYcwF
E/XlZEpDorl+nTz7KvAt59aRY+rEJayCvXmpE4mL1kP3qcPLDvzFLzlskBHm1nyemDViErIlILH2
dYGU2PqwZD6opP8/COimo9iQbhTB8RAv3HEpth1ra0YxPXDxB8F7oC/zOSbIUpxmEYPuXFMHRWD/
c0t1/e+P2M2oM05I1zTscRZrGzxmTu/y5ktJTYi+35IhZt+upbzhSk1vu8b839+zy+30KsdGTn1u
xl/H8AGN0FathM+iGf+vhbbF7nAgSz0ayx80OYH+zMTL+QuUoTJM3HZqTOnvuqXS7XToT7VMWuQH
FTmWgJTM/T53UzznVPAr4s4K4rwRXfl6TMTt/EK748rgA8IJZ/VSE8uc+9OqfQkHn0dfIODUOjQq
k0Qp8GE3vXQ12PRTiXGTu9qYlepf9p5cAiKt0oVAFiXAajnxPqyd45U/53aA/gXdTQpQsPq8JjPF
Tu80moKFO1rHNx88zNrBWgLK40pWDB46adWBTx3zmOa9m7VexKCmX0MNyJmdlj7QVx1tqcgCWJQo
lv2TV9pnih3vHRykhkDej3xa+mzHFpMUHWsWSsIp6sTO/7s5oV6S869Ej2P3E02pn+eYLWjSxvrB
aFSCPx8wfdrfKD8HOWPr+tffeb7Ft8z/5gmA/TBrmub8sASMqgHRFB2u+LVAZjOhy9waszM4j5uD
VN36XDVz0Pb78nv9iQ3BljuZiyPZQfp3drmeh9X80CQgsiQ2sjj/Cdv7wKy9jBFf+ZWsPZdOTMy1
R7vg1dGSJ5nkqMQAMounBvEtLiy3SqQxmiCXhsHTs/WeX/X7YnZUxrlQmuELP4LpEP6FdUZ4IKQ/
0lTmmzabYlNqmTUuMwNN6JHzD/QwcGegHzfTYt4vW+LNuFkdNeCorOSJMRCzCeL+1MuKfM2f//N2
T/24zMKhxvCx/pUkj2GqemNHZA6DCcwDWgfjbKqhjVdi0zyyHomsBG8/FXy+jGcorpMms9X8U5T4
wU2mC9WU2raYaVxTjGua/OU4+Oek8ODpLhI6hN/XjLjrv0MhVqi0+m9uyqMncuewL9ffoEVSpFBD
uxqh1ld3d1A4mLj6e9oW0sUMbgwoz8L88nUD11xIWXkcjreyuKlGB+c4mYF8tVg5bZ7x4oSpWyFK
Wu+0Nk/sDEGWvzZF2oEPfwMnizuhQMIELg/65gejF/JyNfFCjhKDV86gLYUsUXbGtLb7oqF6ChYF
JnC6uTvJzbFAVBZlSsIUu6eC+ufYqRmXwztf4xSmcv4HM72vddWDwtQkZIURpYFO4PAVsDY1aA0p
5ZIfZdEb99vtBid4V4UV6poUAajStrX2MBPnmP0BaGKv73JECw5ElHeFQzh3D+I89094uyOd+DoV
gpcGYZ+fZnb0S0GSbG+KwO5vclvhyxIGgNbk10Z60ttQWkFcIzbKxr9YSxZD7AVxToYfomI7HF2u
kTtsqEM9SqHUJY01NjINXktyoMC+gAY03ZgeXqzNKo83P3UTNZTcuFfc2K2Q/HvyB5QWs9jDUPFQ
Cxwcx209YpWRU0gKrtsu2D4nFP6YXLlMXMP51nHgZhrGEO21JOlLKQs2MQ0CIdNIc/LuD86270Iq
UUMod5O8zwJz0/ggHXIfdtA26/VipbTTJkJfNEzeYEtNETU9Qrfk7fx+LZhIdtbQzet1IQh3cdog
sq3GT9JhHOBwTec9CNCHmAyDtWmas3TJmDa4VxZNw5CTKUhfMkGA/CGu7qMfw3IiJ3bGG3u4mmNE
FKw0CVcPVb/zsNGFmKSPqBmwmrxNAsEfkQbqCjNIGWqtzlkLI8UatvM7o/CTU2QkTtgcnNiae2KV
Y8A0+++qmSHCRUw/XnJQxYyu/NXjwPbwjaIFDirk1J/JJ0Z/ojfaZUM+W6vCTq6WGV9ybxXmL3K/
hrte+fQx6QFklQkzysu1R++19wTCeEI24pCXsojuTDYPmEFfJihJWdD34HZ4AJrSMfIN6br35klD
QvxxBrXbNF135f/desnTZxVUJDMV7q9FBppA6uLHv3VqHD+zi/xDKQ3URWk1pfM3/WZTinkZWxVW
8uFE2pxlef4jveaQo1hNjDnxFws9HdImM3zs3/3jICptK9eNsMz9IVSImuTGHayTFSbS3+RyCP+v
g5yIRfZnJ60Isa95cCjJSV/QXBHXO+PwXYP+rrOMtU7boYwrEYRQGz+VbWFKccr9Ap9uJN03og6U
zqHZC3Ry+D6EoZsLFze6gif0bE0B+9+D94jrkVjWpQre9ZO+lcYl6T9tx5fA9lSc1xlj5uzO157Y
4q9V5x1i5dLXkbCJp73ix90sqUxz9YwSELt7K80BSJzJI8y0AxJfyh3rarxBRK1Go/iUxoBk1BCR
eJtl+JpI+qGmUD2TCJxnop8TdR83UuCJGbUpCOoDcoJPnscFmXx0+LBq93uyautpOIAWBmc+ro7L
fVe8l6iHlHI5ahJCLQgAOKrpE/EmUlqxPlJdJHvbj3x99LWtt5CufmaIToau4CGhgDZNUlpRqhAJ
6PwH0p0TQ2pMo7H3GDTovNzV3WZyNtat1fmrSxuuELgtDm29sXtkt4KCcyE+Yst+zZniQMHuZEz2
ON4kHqubNduOY3vKVQKsUqrt54Bf5I6gIDFlUIbhFUFBOeW43egd5LTQgZRzfmXLi7ssCn8fQn5s
hmPL63lToO1AwoFjUuXX7qr7AcnGx4E0duPuLSUOxpbixDgrndNk9FFsf4AGQXwX4MRdneGzAjMx
yW7+YTHtfV1TP1On/wcmZW4321uyy2IH9GcLXzJuy+dSXRKQZ5uzbz4Rsni431/dAdrWnj1/vFx2
+zD2VQTOamsmphv0zSb2Bff2+J5fLm7wgvvtOsa4oOnnuXbTqWrEw1tJ1IZvnbJ/YI+FRaf8Y8BJ
HUN2SpbU4W6vLeG9U5QyUVoPqk++/wLVOtjxwYdj+9eYsdyAO3yXBSxFniQy3FkH9nf9+/F5vHR9
6id3POY8tZAVnAlo1c+g+IC+Y7LfiYN6KhX5wyRsuW9Qjnip2Wc4DNmn689JfltLnoj+F1eho5i5
5newaLrxTPpssXJJX+3TfQoH2YKaKoOw6rR3DHWDpobW0I1JnNSb1+oX2igzS4cXyuGwbaAvtN/J
p+3bQeEkBwbPVACp5AwCZLIuGyP0vzM/AfTzDf5GTIpfnF2cewXFevoFNMJ7AhHMpn0EuXt/ggNI
LDSL+yGcmXpdCcs3YOVwBedY+SAxTkbiLcf9iYg1Gwe+JGsOHfcANPrDThc3XiIDygGzNiLM+qaR
xKbm1mKsEVTQLxN++b7HGWSf/stXVVzQMX8tU5eDewFcWPprtNWHHn/qaZ/zueFYhPqWZk+biX0E
eDNNU2vQtQLyNIWURgY4sG0It9+B8SD+R6ACguCNZ4I/PaD6ByYNzc0Xt4U1F8qPm2PsS+gAqxbn
ZZ84CntxhF7WD51GnAmD8cpSaWgEWY8PQgZ0vD+mFQyrg0pzdFTqdv3z33PyfwbgKA+uQfSMZHBE
Bv7uQH2fHZl9+FrsTggdG3U2IXujzi3TOVkzvB0ziNpawWVKHjGm9rk8HWJlmaNXUHhTkx0/nMpm
rGCVwD9Nw35Nq9Xp8ZV/UM6/2mLulz2iB2+7Zu6+OI6o3x6+btl9IDnR7ZDnE5hNzJ2Oo2bnmovg
T70FbrRR143mHP4xYg4dxvB7iIjreS1nugNgPQtPaAgYVjSYESz1cCvliUuXlXo1Nl37/fqhyGL+
/XfpqKMKlYI3H7iRRxi53c0LypaSI/UOZwG1FMjueTFMkowiGII3RyZm4tT2makrCVgwyGkLHfkR
ylXUOaveZCxDvZBATj49ox/WyQrPPgCADrC69/1ZHUrvYN7yK65rvvss1DdHdS8naiA7ljzYwXws
mM/pu7SUmQ15MoxhO/iTKwZCeMlp5TCVu17nOXHpdOTHlQdkU0/2IihbNZJIbDIvzvbIF10lT8CI
vuwc4IXXifT0L2vy8XBNyHQmvJcpFbDtKBL9/ekxVK06vUfpfkFczrp65CDsyBWTEzNbrAFc45sL
bsdQaNe1pIFDQbBB4AW2mnEmVGkBn/IhL7IAN2lFHyJJwqohwRqbo3TmjrGZ5FEIuz0uvSO8kVVD
6UOeAfZQz9ZJqEVuycD66pye72dwQCB4RHd7aYRWouPvO+Uu07xYLsnlUDiUJXPLBNR8GseX0j4e
fqo72lqSqczVS1iB+hP5U9vxySNrw9xQQ1LtfUgLkxXU+9Hy2dJSxxn831KgRMiWA/8EYmOgLbLH
wPrjd5HwOaOIqVBu5c/WeJ8ca5v/GRwCvhpHh7954o8DLx7EcnJWlb+zWp+IjPC4Zi7NP4zMWMHg
I5BhK7FzUowyD9EBp7q50A/KiT25Lyr9sbOAcjhjo3dGPff7SxjRukQEDxFyNUs1zQbZRpFeedVj
I9MRzcskT6ara+e/oW+ad8tNzRroUi2ia2JNAdBfj+V9IqtGSEQHYXGlMmAuZ3GBkDUdKwrjbJEB
Ow+JmaoufjWC/9fjjZ/jiVYgLMfb5teSO9i4iQEEFe0Aop8cjPMPNsMdShqJGwoVMgHm3EzBE0sU
/3e63utABm+W27N7Yfn37Px0MHd3U/1bdfi8GFkfMHSuLhLzKk9215APx9AHL2q6HnNuPJt5IO7J
hXM/9lTRKHVqIhhMaMz/YHhvvllp31CmeCetSgXSXzEY9Qnr59fc3LNf2cb1LKGaOcn78qLe0Lds
shwqc2f7ZyZal+b/2y+5/9/+yqd38Ge2b7kUGg/ZbY+hb2jhEe9r/3lHqEzuCNW2ZjKiwOrvueI3
+kk32JbNC9BnH+5UNXSyjJ5uZgd+8Bx7z6DhdUoehY8s2aFxP9mLp4/iN4fs/ZjPjr7kO8ElDap5
Wo4bgnKH43EcwnjxFGagyE6a0CRD/GGbQsMnvlS3t2QQcYzzdqFwaa2gEzXP5X1BFhQR8LN2qvxa
PtdnFGGrUrZYM2r+8eF6boSXMLZJxlFRevLMgz7bfWali7NTYtXgvOIlw+ki31GWGkiuYmFpe5fc
RonDj4MUlwgASTi/zYb43xdWs6R6e+6hOeEqczKXNBrrKA/Y9rACfgg33NsPNNTyqWlV8yvbHOCW
PlH1EXZBQ4dH9h6l6SHcXhSFAQ0aIuAP5E7nqjH1DLZENbKoAuCYFFXmLeitKbPvkhxnL1E+DhAw
6UJXhsRq5yTJl5Iw3zkmnyreodOH/lcfHFte8FX+fgoe+Pdug/DrefDsxHS4Jvd5dGj92ykGWeyv
AKHkOlKDYoyh0MzRMaKW/6Ydfgoy8Hn0+SY7LHTjYKyWaKom8bTA+UwS3qVUpqthbzJF9PQisNf0
KoUi1HpnshhHY6Cv140cEEJyHdjnQg97w7YqMdGir+xLtw/UdTpfgugDUx73u8ToM3ygngf/JMXj
uvD7slHa6Ql9n8Qt1PrefdJsZHzuLbuQf/Je6CDARJiMpETEXph6JTh4fDg356PnkCqIRHEiwHlO
RZa8AjxJCZH0QwKvTXx07D2egrlLKA7tkXFg8tqOVoFxq1n7jsqjJWQMn/RKYNndZdriGzWPD+ED
72mESqssjQYzDkGrT0J0DZLO8vTRq1cYvMnlkF4S9YxwuNKMl5A5MQLYuKkq521TcHqdvHfOtQ69
lJO/OqFONum9i9y09IRPPSpg40AuxBqS/TvaXw7aZ3EaPZixX5L93bOP211cZvK7m1o9z/vseGiq
Rir3Ocgt5ipoGBAZLfRjapWvq8zAhEIp6OV3BZV8gjyix0R0fB8Hj4QZVzRd6iZbYdTixSmnGTHE
Fa8ISM5iO4m0xXUU9ER4Ss8kMStwyRfBnOLlPTB5DAQocFXuszLHobb5lGLKV5EBa92vsKcxstqV
8l/5OlCsV7qs2AMlRX9Fn2uG9hUXd3KY4xzbGUlAEJxQ6PQ5I1AxNPymAPJMb6s9vVV763RIEIqU
qDEYwLemWh6uhPMaRitxSKeX/7/P95/Vg79xq5pxvHhbgd/UCPUWwoz2NB6akIX984K4E3uk/bXp
MmJRuVLlLVVm0VRrHjR82enbfhZoUia2uffCfwcV7XBz0pCiLLA/VdKvUXIgowhRmLKDoNcBCk2c
EcBFZXSQj8pDvmwJ/oEyRIfhrMppgRpN0Lu1HJtLg6sG475st6n0Aooh8UqVLHRqVbIZmGWp5iJT
+SYtU8VEMSeFzYqx1UbxSHqaDmVJcyfPLZMoVCcdb/yi7aniZIury6Rnhojm/xwdvnnPSdHvqfAQ
6elWTh1+YGgTI3Dr4VISFeN/w/dw/L1NY4zsBjeU5ClGY4p0rBGSh4ayrxQP4Q3ihnfYFKiVLrmQ
ylheNg2Eyw2EA1wDVaDC9FTQkBgp95/tG7sEOQYsTVI6rg7C4Ub4xR4UBpP53JWN2gRFOqLCR/+p
jNoRDqFwZ0c8Z3PkyEIlxfgHZmFOfP3jALuPYGEioJVtHRzLZsCM9PZD/MWsYqovOOW/8zSPAXlu
LIlDWb4o8DVW7R/3LPI6EJSb+0yE8cPf09f5kX0SsYxjTtORGNimMZmtbAFPncnKMhLwSnE01aT3
mnP7JQRrGPJ5chVuO1/DfgH4nkowEEJ08TiXec4NroGNa+sfKUycqeWkX3y79JwCzvgTcwHogc+I
vNO3xvBUE3yR2nHwuRvh99+awQtBvD489jRMV643h5+1qVoNWJyBcEGmI6b9GgCAWgqNhhjx+vXA
r1+MrpxwJoaj0n2YWvPq+90Fl62bLb+gJwH1wAtx0yNbvjq1Y3OieNUfAyl22g/hwkb3RIGhvX57
6CA5n0Lc03XIL6/T8gByFEhOI6ZEdlyBUibpIsp6/rG/IXKPvvnGO2X9OUY0TarZKgsJG9fGRCSP
hNl2f+U6CwFLgKugKU2Ia9jjexf8Y/a8llfxt4MKzfW7G9arAIM/ZXrFQ0dpdc+sOgGfwHhOoTK6
/Ch/zjfXGxWWqLCzlSEHg2gJn46CBocnR8VrvTELRj0LpQinGUUgeHWy0y/m1OFsWsMw7w1Oyrjw
R6vwPImTdh1Na39u2D3Ek9J4BfPVtSWNASxpxVWxhKzfbLRqyyW3UWb/iIv+adiVtINwTWxGAx8j
IB+lOnburb5iht1ZXkDoowLnO6utuL5es5QzeEMc8aFXDi1L8OxFNBJxZDd17uVkSRYxfarm32bw
4h2ez7yifhwncr27bmdsviIZsClfdirly5B+D7uKJeMfSedGFy+GcgOLxjN7g7pbjy1DdQYzd7k0
EY431tr6cbWDY4A5HKPPiJMeAmhTjSrPOQO2Y6620QofV3YyoyZZOH7nvROtw3LxofNbBhjrA6EJ
fxA5pkvY1lSGfu+q/i/Rj13CNZS4WxNdLI3+OUrdM37JvqNU44xgjQEk7XJnp1kDAuiixkn7FyXM
EpRpdX1+xl7lz1b+4e9MYB88MwsEWjC8Jy8Eqd6kWzZKM/XMKFXsyHc7ywCaRP6dfAbW0iAiushQ
+fPizXfZTNM2bbmwzPfgnQlJq2nmqaAqrAlMykmzTKIF5C585fith2PVpWbe/ux5AhPlMJcI7v1W
BPHvTl6ReIocvNBLS87x3j8QDf4HXxl+VaMCAWcCzXWAhVihnk/f48gqceOqHKbNvJUZb4YH0DkY
oitFqYMXeCO9O7DT6guNgaTAu5QraxVRfoZ9ZLiRlfmzu4QkMxLAvBUjDDm5D3v2xRuCn/bTkgyi
5N29GzdHqezAsFhzuu/MbzX6mOj9syLd1w2Lx4b+spMl6PouvX5z2VSKTesk7xrMp9H3ABpDADBO
yCm40bdNCLD2XKexPNtBbb2DU2xLuo4dcjH7qEE8iftP5I/0aDFmv6CVSXvoll8hradKtqg/duSx
f4oEuMrOsXVyRlbjIQMy/N/ef0Xku9B9XMBnsppn6ibQt8114cLCBlCtCtkSVSIKRqF0TH41U/+P
G+BF/ahmTu81y7hOovaHK6FrQsrBojbH02ukfXWoaL3YeNQRXJizeC8aMhqR3pqgYLl3j1K8neLC
1v7Ff/HZwHCeFgJ7Nu+3s9HcvXJqeEhBNk/uYDuC6JJ8jOWajDHPiWNKeclJl9bbVpPde2RWhXGj
3NzSA2CLW3Ie0vpUwQbiDijZnivddtEulr2CmNNDYWgsi5Dz72DfTzTWZGBNx30LMwc8wHCd8NAG
RllVKv2Gm3jGlCPgrJ82NKIAz8KXaZ5GndJfc0qucsKfuS2OThniqaxI7bXoQBDpeQhWq58bLSpa
LHjC914yQcDfuTr2auQFS0/WClTsXGDUSN2Mxp6iJ3np85YSpUyLjNTRlOQQ6/158alPxL3a3I0L
iY0mt1j4AXJXGN2qFvA7H5/S6E/qu1T5+LZQu1OJW0zpZed2+ce6RvYWYCfm9tfst5bfxbrQP/WX
OAeoWhOBkCKb6aYq6zz3s5gF4vMNvePyuMiMv9+6qvL2BlxD890omA8is7UMwqjErwQwYmTVVlSg
izJ8bNB8Ri7OII6Si4puf96UG+hifldG2KtRVmennyH/kcTEwji3+osAZhaGzgQ9EpqeEj59QL2h
GGMSJt92TgEhW+xlwxEOs6/teDuSY6F5G9G3ZqRTK192upTsa+c2FeR7pW/M+9AMncvcKUVozDMi
qlyuPtpZQckkpAvi15j0DL8Xs6IBMsfdvbPxH3YRuU/s1rlLORVtT/fl6/fr+l+QOuHeKMER8pgr
Vy4XDMx8ZkPH+e7/6MjdEtieNfxQEL9h24HVxtsJ+DMIIdDy0RJ7FDcGfiTuXLZs2OBbFnKpk/EH
NL/NV5pQitqyuM39xIYRPZLcd0bTICbABtTEV1HBqiRYwIGT7r2B+moJj18aM/LY6glRC9KTdJMr
FEvwtlrHk6UyvjT4toI7AzDhzf2HHQ5qoLdsnOeNdsBN83BbWB0qX7W0YuGUS4/Scpg2diQDEpn/
x/B96qaol5MSai2pIhmKweRarulQVjo1p2Yvj+L+Mj1d2bQD/OSjRBzbPoSJITBMPAW54hiuvC4K
fDqy5l22/xa3NgWljdM2wR1oA8AInBWJwIDGN6zAf5Ks26p6CELd45SW8qgeKBLciHPUtY+yzRai
EaVD7RTTlUYCkYX4ZPLMNN+cZsNWNps1i9F1JD2khkh69r8McI1IxlepPpnQ0M3TsVAfgRx8EgBZ
EaW12wNlyx4sSQ0areMdJna7RqqP0xse0v18Taxn9r7KNzfeRwFF5LRaTlmIrSGJOYCJM510F+VC
D8YHNF2FwHWqqwmxTCTynShX82BRalEdohcU8qzkOrqmNqfrcOin5FT5wbg+OWf31SE5YZDbCWdS
23JhsiLQCh1f453mciv6PJKg6ZU2Or2agqCsRRhi5j2T1Yu77w7HRrib/+ze/erzE1PlE4P4DFP4
TZ4+h6pEQ/BYYIVCE5fPLP4qc9cFcX9K+puC5f9BGg7l0kAJT5YEGhGqK3uJxlNnIIlDYuGFq+tK
TSQIGHV9eP1OVpC4UHvO+PXuEVVh5EAXzzT0T9Yq2NsmbDaPtzjIF2RfEyPfsbSXy+QcLDsdVhPP
jSnNiSQkIcPZ4savk1j4Jo2vsrwU8OmMgc1oG6UodAoAn8mbj0kEJ5SN9Smxj0GIpbmXHl8wxffK
tra49GDFrfxlloXn9jxK+rXP70f6A9WmGjKE8WP2R401ZmXL8AAGCmVRCtN4q0vE3SAad1uH0fc4
ScwW+jHT+sJEQe9X3cIl4j2wzkEMl6b+Ylq80p5yjbzsFzxf09WAxzKwk467Ht8A2lVSlL3wZ3Za
Cv2tBca3DHMiD6wRRJg6vtNp/KICjTEiY3TWkrIHzohxPeh2JyThytdLww9jOQU8zGx6FAB7bkFJ
p5P0r+YdVduMySDnjPb6ZF011zY35PD0Bkchj9Mmo6klYT5Od39viHTu98dZPy0kGKm3WSfRBMu3
v0O+Y7MEmaCjtqYdNFqLygpHbI6ZowWPF9l0ka8llrb0oKHztUGNCnnMaY+IEmQYj8QxOWsxxYn1
aZcUvP5T31woLxvu4/uRiOlA7l6hmJFsmWCJNji/yJVzqQmWorv9Q4Di6OUxporHwV4tblsxm1sh
pq/6HhaBlHUk7wgNqjKPSj//u50ZKPtiBt7kWpjVzH0mw/myVpsqM8/jVXYenfpTBptgFQBvLu5d
EMV662G22hA26xaiSk11h7TXBt475jc/mg4FZuIqBwwyO7zUkIxWSAbW2GDPE7qEnMlf6lGnNtIy
ZJjwz9TzF2eaHZKYtyMIk4I/Kt7UMn/OoL5ss2RtanzmUXr0WuuWTO8aa6qppQj60maX63Ov/oEF
7KNCKI8YgDQnbtcKZH7df2CY1Or1Tuxs2cmQxmwx6G7+y06pWWh+5NnvNxgxQwzqOKnnIUanex+J
BAzJf1oAvTDeRLshAAyuXIgn447qkesJ6vtrPIzV+65oYJPNHyWyWaXGKCUYsfEedWcWBP+TPGqZ
7e2voxgOIfdlCKf/Kdf2GDcSch6pI4NZ4Sioj0lGnYPzMiChzSW3y8ayg4igGMkrOu0hbtN9YXVL
XxEE033Lk7+ZtweZZV8XfB90qgVdAgFeSeyBgR5H+fCEWEoujXfr3j0S63P5fwd7TQwD1oeK2ZvT
x9zCuw0UAQV0czqrfwvekl8uT1dP5z58cDqM1Ft4VUW83CoXtv8XQzueamUsnX/aYJetkmJwJALu
vzqiJHR58cJ47V8im3/GSPJV+hjBY3tlYSENa9Tg1eHNpMPTF10E1oEKZ5lOPIkQVMI2GpaCXHu3
oRvo+w0uqXSsGvtPJIdVAkFFkViaZ4HxNRQPrFVzcS44wPjlBPxRl+vhpbgOWal9vPKU4CGNxkxz
RsEj0/vwk9M12v4HwLwdcx/wcBdJrrq+NNaImmihQdwnI3F3oOM7vTMOAzqvj0f0sFjcwgVcSfhm
RL1FdVy/oUxaOC3h1ATcT3vvYXnF2mVgs4nsEBlTJO9p3f+Z/vfLHkxEobCDt+Y+3wDkZ6VWf8oB
KzyVQGyYTKtfMDoDc4beAgaRDYRLa5QrAkSSbaLgSGjp21pER70ODAcFnzLE84+ASEg06Utylg0I
2XnzsibLn6OV0ntnRm7NfuFdtKjqH0svPZkic6OVVNxIsWP7ZPGDJGNrUV+Ut/KIfICAzsYEshGu
agP56FaQil2BcKZIIfB+Ivu2k/Np1quMfmUHg3RAiBpGPjKBFgq1NvefQ2c0VRIo5sY1iLTNoPLh
lglmyK5A5TKJ+ilVYtrDlSoh4roemur+s58EJ7+1Uuniwj2GnDljcRuoMVifVBn7kV+/WwPKFqKP
kpifEetRLfHlMCzZ/HXm2PZaAyFmX1ws0vi4Z5Bjvr+yC++7odEVtbnTc8fTA+A4Rv2iSqWZfN61
QMRck3QplZYhGcTbXvEOGlF/thKzNp/+WOIu7bEpKUJ0QrAySLYTQkHxuKfFzVtyPnv9w0D18ZHa
DNXNbSY24MH22VH21Si9r2GLHZh323fGUryH8jjrzAHky6JidjPNbfBifke0uRU0vsNI5niAZSB+
0eY23lB482RuwdPaVwhdovf9080HbyTRERGUER6xbjWiHkPw6KgCxSxLyghyj3U9bQENQy9onr9E
9H3pFj2364A6CklCQUmnxh29iS17YeiCRU+oTQSj3XN7pF9waDZJoEkY1vSJ8kkcgEdW5EKCVC+G
ChQkCAbSMxuoKAdJhAv8aKcxDUKR+XFvWoZYRZW0Xb0F0QIxP5ztL3Bs6gHkT+qIaECrhpMAFNN2
zCFXrjS4A4GT8CfWcB0Z96nbsSGqs1LAMVrTiNUkEcjuzvtmstUkphQle5WrxQc+DKggmFKfn5zb
nLw7J9Kj8MHwwYQ6HKcdOQ2bHayHFkyUMxtkrosaBlSymtDJH0ddTRTyeW5Xl2zjB3MzcERFX+NM
Bl6pJ8xFm/48trJj8PjdlpO7zHBQ7cnJZcpsGGh/wg84synw1bPi7BYXZKJ304Nk4Vz9/Z3SFhOB
G8GWK/8sHC9bMdOclg2BAZhuFxo0yMS0QN3HnHTXgPev3DHp/aEDUk/bRJW8Tz3DhNcXfcUfuR2d
iAhIcBKowS1QaTpbQP7i6I3dv2Mhr3L9SzCbtd0K7Bt6Ese0d8iQuYP/Q8huNPGAJHNnbsQU1qIg
uL/B9/d2P3Aw9UDTE6fxJtv90jKxeiMIIJqLQVQo+rtoqIbMFqzPC+2pTewGn/9JfLQ+6dPbQ3YJ
Zzy3ZoYPv52pjZI8LotmAgnP78u3+9DWEOzhy7XucQttZ6seNpamnNzd67R7N37d2/yl+rYPxAfp
ip3SO23W7P4kMLbQW8Zffks8t7erH/yMKVz7dc642UCHueui6yx+mybR2pqvNtoedPvJ3i+8+2bP
Qg6Fw4e/N1z0Z2ZGOTM5aNCuXshXAs37/cZV45/T5q/ZjJ5UqK43ObCq3DvBK3vHk8RmK/1O87iB
QTpiBgcgK1ER9HMOGjSjlQqNYYtdFmjnsGJoLVh+bYvWi3M0EbGIjGQCLq44Wcrp9SAc/aA7p+Jk
dRfghhazXIONDsNGxGtprqaV3pRHAzGpLCUDUFi0JVKr3rKEC1maS+DfmzFtksUC/Pmzsr/vssMf
X26ce+iHTqj/5JbcuV02+3s7q3aEfmuRPdeOlXYOLsQ6aAQkG2yHq9Aj7WL9xVbOnxXLk95IRxyf
qqxzb+yQtgpcyD6m7YtkaKCwkeuxPlkcVb70o3M7jycNmyYlLQ4huSQFeLZjk/ZQePPiAArVbLa4
N+P3jDj9ssYa+n88F6uySabCig285oSEQs4rgdNKTmblM4IVWCJnH9MNsoLO/Dna/WY1ETRDXfsQ
DbHx8Cb2RWDAQxyEC0JKTahyJipO4nKDs+7vg5ssPx6Tn2g8wZnJSTEIzqOsfe0AgVZSli5TSCSQ
JM8wJLRaJgRtB+b7jjG5Kl8qET1zYPtZ9S8yj11bWzcZ18yG6wVzfnPhLRNwOmoj6u8gcUqpt/Ch
7ka9hxkNMi6QIHsQucnGXCbiql6ufhHe0zgGsn99KN6FY2otcUvhnh8BY0O87mPsGf6KNko9Ld6n
IDRPUVW2T/u8Dn0f7y9m0SVXhBr5elxISUPODZsUrg2eBFlIfLgQxZK6plb2h8UMviJJdgIsBsfJ
aiHFg1yXPyDP9wQXLsdIl05vUKnIAMqvdDnlPn6cR0SV+vcKETFW8WGsueZZdMS7YPuKOu3Rczdf
D07tO8j+OmcPzjqjpITgqhzTAmmHacdKeehE+VRq+S31ZdkwVvgONVB7lJnGPMAPSAqwo3SuR6/Z
oCrhP/oQ5tZZlMLiXHAhIePBdZBpxM3zCmKIPbENfml1uA32z6qB4xkAoG4PlTjfAZdr3yekgGGo
h45etzM7yhR5nt/dFoEwelWw+jpbdCCcFG1nTKy1dMoMhwHYH6quJi6i4lInCxZaKd4Kiu50ka0N
sZw+sTxe/n311J1NIyV4U0T3iWG2wrnoAS+OGb18RlGO9mwM4O5dwWbvzbrRNUreCTqIDEeHOlW6
XiqSGiQmb/NLw6vaKQUry/dCoosqPrZJAGO+SH3+/08acsNoFb/C9MWk40oWTq6/fPG2IYPqTyUa
cbunIe3N9we4UJ0mYKKQyB8RlXcBmEjjAyHs1LwcsaEQHtkNc13loekcLmNwY0yq3tZ7yDaGy6NY
Ec+mivhJ/dhI0n8um7Mfk/DVKA0tMY7ZXYvuW9yI8YizZgjbHPqnZf7qGtPw3KHMs7U4+X2DAJOy
5JtpZwn+huXGZYAdtM1xb+2ZTcJJ2phtLTKk14DRYvKLV7dYp1mXmO+dvi1J9iBW5aL3eJpH6bol
x6PhzG3nroXNwtcViNLrPrXXTQXGdf6e7QRK19lccVhLBEvM7i4O28n5O5NNK0SkbAmHDdIZ8F9I
GtFcN50thVk1m39ZqocjLpETcM9IuisbRKTecJ457PwMKjwd5hmcjm56Rw5r+gVXVZqMMWx9xVyZ
xKWt2oA8EQcJ1j8+xurZLp72FdGNONE40A4vFMlxv6hUhp3lq2K4v0yxmO2jW7pImQfiyJaqMm8y
Y6p/Vt457XQXAAw5phO5K2tNda8yothzUncz54r7wyMCMaQbrWfKau8mUdmV6vAc/8CgS+5kmaNE
5YOuIVv0IkRhRTP45nczccRFPOX6yObqRQBXkaEXdfmMhOoj7iOwgz5S3+YysA2ac8YOGvWPSc+q
/LBgPmHo6QYyqKlb4vQbORoigZQagfStoIFoxrubhv8Hd2jA6wrcw64HCOQ5In0HwqXLU2oXwZeG
Stqq0QVC4BHrJLYCI2NBwJfPbUok8QpY8VMMU0j5M/LGSYYyUtE68X7276M3ijvtXINJgxyADgeT
ncuUZXcyIz9rl9Tw2xFMTLOANZyVT5r6DWTAjbj/Rd7x2ZX7jQGmIFH08LjU8pgZAJ9QP4B8hJm+
jmV5HXYWV5T82OJoraUSu/r38sOoolna9Cd4H9W4r5rYmwJgAV9O449OFO6Yz0vZjitoQzag7vik
JfYDLwx58PnfK2uNBDuugvi1PHHaBpOQsg+diT1hJ7LjZA8i+aAIYRc8+JRcG3P5FbTDB9edbIe2
qu1EAq2zwWDyAw8RSJGCU1GM85SAxyCZxsm3pOQ4Nl+yMlCfMARReK6yCPnOPFuTx8Y1Dbr1+6fP
7Kju7FnPUrZDlC9K1+PzE9qW6fpu7G9gdmw47uiY1BSjEef2YqllHuC4wBug0zDanMFL/PeVZw52
w/0zZxieQ+9EBVHb9iQtzADkfbTOKW9Qx8lGKPJMGglyPaOt5Zh6F4addQrrK5VJFAfvyK+xJzBH
fj3ZPk0nVLDTx+ZAGaBEmSmWDp5QizopsUVz+PZmLsEUrocSZ85/cb3aOdvq9gmcVsNkqc8G0gFe
SVuZx6g80/dE01Ur0R3b0tPKAj29CrwxZkRo0/UbNUxWz6QV1kz2C6ShI5s2ntYkWHdp3H+qGW/9
BfWeKi6CYazW67zK4guEWWYvZFOzyYFULYZf+Uhm+XRdtBYgIxP4bMh2A8Y4PTZiIocrWmhZw/KU
H7FgHJaaC/TtV3ou00DHYQoHoZR6teJjQXyw4m01ePvG8cCE7CpohXoapY/uJZod2jzmrSlYdBgD
foNJ9a20oI2cz0eqIJ54zG3zrDRpG9oIVjbTOAofkyp9bWM/eM+pp3Z9xMXdO+qCCarzD2WPuTZR
zW0AYJxo/vkTf+Fum9iGcwx0a7HwwjWDY8+R/+X7ajpTpoUNNMN6duhpgWuUUWUgjgrGpJ6/j9Eg
9f6m6lXZ11sz6+EFZFlg48mRzAlWNz7aHfQJACO7i1K99adn74r/qYwA+GB33AzOcSXw3UlS1/jf
zWsubhfu5+LRZZFF4gmjBDCWrVTcFxA3Z40AH6tiD2xUQltgzkyB8UfXhjKnvTABYxTk97vHxfrC
NQwGGMpnnfVgqYpuk9hzmZ2wNb9m9fKpx787ojSGWfcvL2laxzjz05CEun5HPnNTHsFzegUWVi09
FbQYXaJbgV8hHeKhhrOtvhjL/QhYAjiS+o9kIXLuUO/VPaAflK8Icl4RNf1gZVXWyn+WqrJmfl2b
Knjg1sbFm+py9ooKRm0sB8p0wETb6PTWjzekcl3XQ+ymfZ5wFHvB/YHa7kFDnQ0Ys7trYd9HYaCB
b48rjLwQ64tUUFWGfgH6ibvAe4ypfjmOybXkv5ZoBYOAMKdtNg3B6/4NiVP+1SqQijCqBjJyM1BO
CKU+pdV7WHcJ375xXMY4FRK3Rmslwykp2YV6kLw/aBNCpl9ABIw3Qn1mbmdkC84WF0DjMLn2CjQi
VT80gWZeH4lfhUnZ9Ew+KUw3HQ3Fe+6u0Q4ePLHyDoFyQ18kHeD7MgtOGDA4sTBEZ3SLYUjUjQC8
nc35quj6JCrqSKTfMT+ZwaiPx+MGY+Xz9E6ITejXyiYo9NePXjSQGneI4XoGHuaS84Q+caen59Gu
7Re1WI1phVNeeALnteWV80eIP9Cq3DsOH2lKkNHsVRKtjkrzP6DHtfVbTq6xwtjE6lP5qS6iWi3g
h1I1SiKyH2Pz33DWqktp9Ln5wlaqyvCEkBz1xLO9kVNwKxwbtfllu4BThMtot8DUB9US7Avl2F6I
FQdZoHSTTkhkewClr/ZKsXgQ6WmkQTmYdGAusaytpRlCA/paeJ5l0+bjhescV2eHyFTjm6CsaIuM
1TGNDDGimsBR3i3Ubu86NsaF4pxZX3WiwyuPfdaHzp9cAlfBRACDcQzE0pb5W8a6mD3zI2v+EV60
Qr4Mf4vmgau1KYFqdLlQp1aMJM/R+8vBT/2P25zKEZnQ/EUapxcRwWbTFcNCb+F9ble+PniRDx6A
2esTGF2kgPWoq4A5cLJx8+IVYDJkNSPrwnejR6BV0nwXsnbBxXTxAhSuTB24ss1InOGYsCbeg4De
ZPZfXnH/zfvjY/MoFsdA0geQl4V4sR0LaNec1TmxlgoAhVRsRJBGWCnn8b1cN9bv1NsFVEkIy9Oy
sABZw6nQMC3JhMuTQyUTkX8UIsLMz/mL4ZIxcjGNjRD+xJ2sgxGQyzj56RR9N4UbGQjnd8/Jz5V+
3x1r4+ytKcLMzDZ3F79326/Sw9v22qlsE0wOc60c8gmhhYKu6jVNPDvJ2UByhnFJRrcxCocShuuX
vwHHokc9UdVEVKlN9TdbmS5WyJ1xJC8U3UxoOJLbR1re1DNf2L9q5Mmk29Bo/yrxuAB9m+EpKIH8
9uKffvaEKvgTDYMHraegFI2za/QHkhvoDCU1VA6nqRa32WqvMVYT00CmVOvLi0zRfPSyJ1F2ziO9
vY+hUPP+RfiBvaflnM9EVaVlIXQzMlkvjLKDPdJioXc7uq33L3aa2Ei5TWTtgsfsRbLK9ApWOqez
X1z7erdUuMawD35YBKSoHLPJ9Fdvc0l4f+uq8wFcztUNOMhpxjGfNDbAKjDijym37c/ojc46lBsT
HSeGv5Z4k74W6dpTFAIO0beenpOqTgWvh43SzQin2FZ/skYVS8FnaJIjEQGTIw3Zca2fOv5khtAH
QvpsA29Ev3yc/CSwf1fv+219ZhQ19TZ3hbxQXp44e554BRwVTTAwLRDqcYiMMtu8WI3AtmJ9H0F1
tYitdmUPrYhIvPHLmANIehJVgc6MHa33+ErJ9KgW2IAi0iqgFxw0/D/cL7TdUUjDMDeovg2sRK8E
vsrRO1r1QsXBxlN1vyEWkDBm0llk7l1OuiObPzmXXtmtmzAmByAJSFhWSr1FuTSSXAfbahHgar1K
c3KJaqVOAo+a3gc9cBPjBlMsdub+luBZeLkDhdTgwzPZPYJ7pNzF/zY5SUYPpp59e0nl9ddzOETH
IzTFRdZ4W1pXEzDVlU3N71FK+RNwLK6HULu7A4yJsXLl2UDcLvgJyYZ2JHhDwAIvIK05IdjsE4Z7
5dUtukMtzqlXsO4L1V8x+z7N/cXe7q+ys48tOA7TSe9E5BCF046k/dhcXLYq6WYWOuvtMDycgqdi
882VLMXEI+EkX9Lh+lqeIB6HPIXg2K1fI+TfcG3sZnTy744IS8kWLaiJx4Iv/mcNXRooiIkJSRDg
Vs+QfG513WwHYRkK6NUgiABnc5kbjw6yGH4m22N+7x7LHD1UXCBgPaPkMTv+543uLS0xFgkGHGf0
IRrjYHnfYllTX15z5j8nh2FDyulOP7prtx/ZFf9tUvZXDed6KbAwfaT8DeW+J7U7I+esCH7NLxUX
K0pWacODVhalfiqJzAUcNmK5aa8eDSM9nPasbyxIsbbAoMG9n5H39NP+6XgEAm5i2Q/Z/rlyOJGZ
5mreUYLrliH3TCqqZvEM1WgEvj/SmUddBVTNqTMaH6+rKbv2+/ZGbuP+SGMBAzJGgNhuxN/ZDhYO
nsK6XfVanIQ424lCvjVs64YhoS11x11UruvgcEnkkHIdLEGRliEnCKknLq2nShS8VpGSwGreSZIJ
t+z/jvFYdTBbrQ6zIsZtKUTXnXTbCYMwh6EDr1mXDWeEs3qE0b0rgF9ybW60fXjjrGwhTtEf+U1G
o2FifoF7WdABwegSkTvAVGSJC7QGdCAe0vmDcy8YRtPKh+pgqPJ7U8oj5d6hKutlu9ellv+0VCyo
77GeJSCe2gPdAWxjfNfHzTKb55VmvNlUTAzjNDSEhB01DiowA7912KEUpUS7WIWGH24fsfpmqHaj
cPqxmI8mdYWT/NffiTI3KmLNmAzWwOX+9p1lR0A8n8kNz+9h5dFiDrPEiUw0kGa98hE2MSw0m96J
JY+NgO6qw7L71h5wOo1VF174u3lUNVwtsaTX0i+mFvaJwBAiLZuN3/hHQN09+o45PXIQ1iT+WiQM
zsXOBbEmL06PtR446oSG3moncz37TpdCDrKsVYlTDqhCPMgudJxVYqC5b6vh+p4IRvDclsOUM5Xq
BGRDJuskxFx1JdcRGgowCYLxo5+BJHip6Kqq7u3x6TEjJhqoJyHTDRbNuDCN+TiAbxZdCS59DSQ7
oAXjPu8pTPEViLq3xdyU+eTFWJuZOGpCxizuQVhiE5fTx/0G5qIrOesnaX0T3wZV/RZRuFPBBjcr
0MsLd1W6vXtBA6gSB2euFWi1ulcmqbhamUV8Kd5OGbKHdsP02+kGo26u+V4f/K0mGABpym8kC9UJ
iW+twjmJLIB6dYv0jBcUG2XoJh+xpr6vOs8tWpuVSmkFXAcMyaN9drL0t1ALxTeem/M8RavL2Q96
nEkjY3I/AeN8wHz3D8sbrE0cYoA16nYVcw7UE2GUwB3LZVFHM2IsF8uBWwB5MEnQshzjXRa6VIJG
Ua45g0HJW3ydq/S1pMgJ2hCkY+C9woFkQsnNElkPB+riCsY8oHa6LjFtQM5RRt4Pd/v7uY0m1pyw
rgooTQyzej3U6VqtXQMP0fp+o9qTLo5zV4T15+rcesb6XvDvTGaL0KGN51vJFgITsc1Q/5EQD+mW
R4TsAyizfDDw4YyDa6U40uc5EqF3jP7RZkpXxpdr3pcGJOk6YYfYI/U09IuFXULIF0Lf11o2tbDU
TdysEF/hp/hHWKR+f0o+ZH/eAPKr+pLINZe5h9+qKt3WZLIfa4vPX/AEsk34zHNpWfnOdMnKZ9oL
sXPXUIrWojN5Y6W+y6kUFIx86F8X7jeoihyHb/96A+k+1WgV0wSD1UayZIXchubTdqPxkwkKQMk=
`protect end_protected
