`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cuwI0oQvU2rXdvYd8Vd+R2ZFV2YLvapLX5K+eUcvPkaPZlSWNYljhoKUMsk1rF8KPQ0n3oqY/PmR
APQSrlrN5g==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jT+OJC+6drO9SSjBZNMePQ6A/gZBokUiLux26Ww+6BdgvQTdxThFIShYudl/QaqAIcXBtncVl2p0
a3w4skbOgFkuajoQRqyt8nmAbRw2Lq54hGsmZ4GYFZF+iQt4UnwkQ2RDm0f84MgJo3Qw2LYTX7mW
o6wZJznKuElYgio3qjs=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VeFZKyTBwCxiTC5U0t8yEANXr2G1x5rtFHR9sBY/DkjWmXYtphV8vQnRfjTkippiM6CThr7d3icX
MPLkQ0bE5aksd7+ho5m1i9HXs3/OQ76W3XTmtCTSiaqZ5k4O6zb2hgoO316D6g4GFfCRDdRSpfn+
+pnM26jRqOFdhZ74pLk7bvkxT92wBogEApg2StHt/ISH3rCSDW2IRoazBLlfBNHBt3xyZawvQHpI
TQAt/G+hRpYHnzanPJbS9j0lhs9PVkPIO1bRO2ndUjlGk33KIJtoLmBg9MvIMwSgKMfd1D8XgG2W
okXXfhnnki926D2cklg9rK3C9vv4IDLh4gkgZw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dQHjUodM4rYEXa0SPzad1IOPsv0vFU5zU3gHQEnVcGHQ5Q7uMimCRjM215XbaDv5qn+Z4RQ+kJoN
HXDsTitMW/D5EYpF+oQMe13HpEhkioLB5LP9OU6/4GkZiPV4egJJPzmWdSXpV1fqnAbdWhYrvrXZ
cUGuLibi3EsbLUVfo+Bx1h+d4EArgRT2G7qJw1ovfMrV3ZWBi5rj0odzF5la7cg2Rh5em2E/lRIp
l4+UwnoZm4Ewo5rWH4J7byZbIEXpAYinzgTvZlGyCScGiH8seCF1L/YTApmJG8gc9pLcCYhujeCf
RXPgKWaIZFGJStq8N3gtLRLxOkDRRRiLo46Ksg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mLO/iEW9mG0NqqzUCPoV6fRdFNsS3CQN71o7tUo0hjHab+TkFpOicx5ldF7bVDUYhynof69fWLUZ
tLG5tIWYL0vegV+AlToC7Z0gnL8oNHZMUt0Aq8Zmo2XybwiNzTi06lMB8ze94vh7c6T54pMcbQGx
nhmdA/+nG8I04ONN2n93naHKp1UkQzUWE7WoFSTySWzWK3CmjYFd0KoB7JxZO0Sj6WGa4FrBwiT6
9OhQfYhqLJTqQbYR2PztML9hchY3qnI1zDrc9UfWatGS/wre0dNE0td7cvtmBCNfbHzLO1YBIdCl
VikRIWca0nanK+VSLuGnNZ2msAlsXVsbfRPefg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
deQzHeQZeVYc0PbXNWoNQBYhCkeUEE0qcOF/6mj5m/eoFV2b/W/YIp39Hc4Pze1/PAkNJTg97W3l
QEJ81Q5bGpJg35rKg5osGcnFyVnE/f9HfGn4sZgdoZ85GgtSnFN0kjzooGpYHmISQQawmMvZ3m+T
NDcU0+118elNPM9uj7s=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
U3noW5d/YgF+qYOMT0ftwT6uLymMsWtKAJ+tEVeXvlFRPOhWjebKw8x3deP0EvN6ERFSp1y/25jg
omPOlScJbhl/biGeTI5yYptBi2OWWGbgVTWBAZl1azjtgeLmZuO06f8avHM0VSNXa0C/IPlivlrx
iof4WpucY2z7g28XjxyVzViD1zKiqv66z8aiDShis12gMuPuO/Zn0riAILM6i0xVMOOWYGtiqshv
uh48qYTzxOFXHcF8GI2sCtzEX2H0JGB8Chxbj9PFoq2JRIEUDqMRNfbCvtbJv1BHPdQGaRHtqdPO
HCVjpOcj1MFbHzC2mzLejxNaZ7Fv81O7pE/iTg==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hiFobri6ZKHb3WS0/M30Yq+e2I/w6f4Kj9htX27P1B1d0J3Oycn1ZDZA6xq4ewLXF+6mYd+yKMS1
mwmib8O8dhRbg699FCT+wYr+ZngDMps4PZhmPbFZ/EPpyeV7tevqB4VaM0jLwzr9UaFPXpCk3qVM
710LUg2B/TIbYiDiHDKfezFs/gZAvgZ+dmMJtt/G8zw2ADfgp/4/P3013IJtOH68HYbWMccCOnlO
FHMKRZix2JgiKMEoho7zV5JikgZM355JW9yp8ZvDoAx8BhGzC10P9f0K36XM6sTxKOvOpRR7ZZYq
tDTyKHngdtm2bk0cebxtEeyddbwWuwMhc38e1w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 71392)
`protect data_block
Um3zZE/zK/gqndbi6L4SPkVDvr/6xdw5EUT1Me8dVCyPLnIa8f29xoaymRrTPnAzjpj7DtZ+kgYh
L8/5ob81LsJUyh8fjz6hi5Gqi+BAt1iEafnGG1xO4uyheV/dIoAXizvybHP8cBdgV4FhCukOwobg
2ASPGyppLvxo/0qoCkAUaD7oLL7s8tZPRrjKGSvj4Vx1Kfcab3h9QP59VjDqHBx6jhfbDW1eJ8J5
8dXSRrS0YSsguk4E+xwb7NrkPW8+D7mqcQu62Rmv30nP00FhZ/5YbvtFUZqY14r4rhr4jjbuaXah
zAqIxs/msr1UZJ4vu4HFjXj6S91HMeHIzqtITx1Xec/jJSxHppbYX0JUHrFR81UufgdGEw0AAv6k
CTNokk+dxt5mvUaqBmwy93sYbzVSTkDklzX0LqVw1fW02ljSu5/zmqtM0ZYyCRDYZ26G305Lwoo3
lg8ApS8tU1fNtEynYPLd+qqjL/bgni0LCSEOmp4b9r/xB1WP4H8I0WRXYMMwDEHROvpfea9A/MOi
qvg5yv2OZ9g6PLcVgKH+SBHD/uurpsi/L5YloKOYdIrd0g6WxBGQtZ5ydkgC7vNzP0vjt1FzuKlZ
GKGmKM2+TCyOvjzwZ7qVsB++3xBU50AjMoEJp5KptegO7PBDFnjeuTm+7lWhHddAUWfax99GeAkg
kdBVhCEOEFw1x9bS8kV7rjxFcXNYpCdMmi0xq2n/QWW7tUMt18LUdlpWouMX3LfugTyuhODaP0v1
T7HLVz3DcGYXHdf9BcPxI3At6PYcacD1IaAfbt/ovXG0RLFNbzzxV5UfJ1eVFErDObRm3I48kHkW
fLCRxm9CIU8LdTlPSMUzbckf6zFJ2/AgM7IkqOG7RGKhu15wkVnHfEIEjSEqXYz+ay95iZQF4D/J
z0Fd7GQUFE12f6qq7hiKrIaJTVyXt+eMqnnNYs+EsxXP/uNKt4s8UwaYIG43S9tyIECH+DGyv3T6
7BpgHyJq1XFWXB4ut44BSxLyTcbW2F5cc5cuRfXHDu2sukYytH92gbj77BBubRgvqgc5PCJRNgAQ
FEPoDh9FzxITG3rkIlUY38qXt6e9A94eJHxoBcF8+/TgTo18MtxV6yeqZdMgVu0mS1mxacLbwRNw
Tq6P5POVC6BdABhfAxxoes8NuQlY9xAidNFCQM5b1QohMF+dk47Fv4QLBJXDAhXFwcWfh8BCdX+z
Zh9xaCriNEI28Zfy5uYjvKNbeqQ//eMExp8R/SxdookuTbHpUyJl6k8ConCkyGOtgdOg3Yd1hyTJ
huJkKKS5eV9KlNdJuWXq3UbuMGWq/GbG5B/Y8Khs7eW5VbPCeY91+v0I53MKfz41wU82gSt8L3kA
LBcwR7gkms35z49tnQirCJVz0fDajrbfysTNYV/b0NnfkRg8UDZ4CHih7Wa5xaU/2nOT9Cw2Wmbu
ABNWtV/JLhKlVNZhpNLqYwU633ZudQtsRUhlUCOTuf1L7BlrVF3KZAVYexKnEznXJM8PHwRoGeZl
7fVbN5x1oEek0wiK2ARqN0rKlcoOl8uYo8Fe2JIAiAd1pZnBPCMbiaaBATo5qHoSJFtcwzDjx1aT
0yA2ShkYimIXziLVN5jOemJrLaTGcSxr9zn/c0/M8J5dUWsxtSnlcFRJT/XnxZvOLUw5+ibKguha
2je0kerxQPgbD4hFScQq6JsAkWd+qVeC8uZM+gJtjrmTNS0Ecxn/Si1Mgz1Pba5u4upz1eHtr5W+
i66nJUPymdd0UDNaAn1H9H3tHQuYKnpQfiOe8TZ+vm6uNb4qKUViPbC+UHGNHZO+zcL4lmFBRdgQ
BDuZ7TC8d9ZrLEmk6ZzdUtNqMNNcssOezjUgQ7+jsmdyHormztU9j8Je8wAJhyKJv/x7GXlNuM1G
zs7s5Qy8KZDmlKJ6WaKpHORKi22gOZysjMsr0fLVQvpq5QHQHuLzR05Y/ALGbyeQo68MijamqV8e
sgbfIyR37zCfYmhxHIEo5A7bUMbJKce2WdZWwBwIRLvBsKF5s56uAgldi0zoDmtK1m41FD9/hHKx
YZEj8krMrDvu1M3/3xb12cFsY5u4MNYLSRWYD/ItBTBZVukfcc8IL6arFaURHed2OFyNUY3MRLmW
uqGsDLwL/PiqCVj7ITa1FQigrYYwbYZEaJgGbUtULFSOcImecZcMKn4ikSidux1i0L3qfxB8kJvW
zRiQzM2ViCRXTHKMNLmDQxO/1Zal6JeJykSPUz7cV0i9WPvOPSsDePZlk/amVkc+sA/5YyjsP+Gt
/pPH4LmVVRzgD8jQl8d++s68tcDXwZYvbnt0hNuOCLjymGoZJa99FxfJkGRcIwIax8Y2vhDwe/6W
zCPwTuowcJAA4rZANOLgVUUUcod8nLdVvpxNThWuCsVY9gEVjYs38JezJx25+/cAVy8VR8g2Ox6O
yj15tIT5wyQj/kcZigGV1AfSgZgTxwBVB8sWy9hBhLEwIYLVNIFizY59JsMtSBQvZpHK2LRahEwD
O6FjJBjIGYIMU4Ff+nvN6Iegt25nArfdd8vWWjIRXmi58z/UxTtfZsKXefO15RU9CfK/3ogPODR6
w1dJn0xRSefPQamouJgSzuZKN35IHpzmlnm5MOjAvaqYlmhlRnyi6WIwz1dK3a0EcVKYdziux3YN
ZStGBXXtmFkNZ/hsD5eUE5Ni1OiwtdY1pTPAglD7Lm2r7R/eMRhr+q+mtS7PoIXde/wyYakzt0v9
q675akfmaBn9bMMElxUd7f8QGqi7h/G0bUEow4dPolb+hnIXXiTjpRyEL+RQJjJn68IYEeAPDIJb
5xdGh8t1JK+UooFLtKy9nzJbwyxJyUUDlERwOvZj/deoORJiTefwVwAqTui6Ww72tYJfJx3ErzyY
6qDCn7VUhtGeU15vn1adAJzChwWo7frh6iSJHuf6pp994vpY2tA6jOhvzAcPi2gbkDT1g0ga0SmP
5ftWF5midWP4ScbkHUer+t6C6w7whnlXNuna2vO0FOB149Y53gcnXXShCbLVruQEnUCcTGRMBnBY
tWvZ2FasdvgoPJbsFyOT8EZ1F8s8sX0/I/quH2Vb6RU7j4yE78f9MOVatTDMvYAheM91v+qo39LP
NjTlT4VcFqs1OehgOFQzNEV7nas/B31Kigsndihn/1BhEwAejt2O0eHBysKl+Tps9yrWwZLKp4kw
C3Oyhboz3plSvpETYT1qQpQbpwaflYdZm+f+q2gofE0NHLca6XQ7E2z0+inv66Ts7u45aeoUBu9j
X2AXBAy5+RjCapA8J9IqkSoi0Q7Q6HFS3YouhzKRcUfGMh8BoDxR1yGQ5VF0p5/O2jHvq39iakaq
1lnh/OwBmhwNeKPeCNjqbl+6ory0sDwV3XHqHBmkF04G8mqbBdufIzJQ3+T4/VflCpO3brnBJ9uK
OPk8T3DA1uEh/Ii7dw4K0JZv2ebJSm46gF65k6ZCiwWeomoDf7x0wVHvu/ot0emCAXi8pOVxcQgm
717YdjhxztM2jCweBUQ4pXRZI/iPTslynrJmjiBEn2DsihQx5h6BoN70+DYetsTJqlZWNO9l6MU7
BET4zOivjeTMeiA7RsdKXfpDv5+eCxRTQS3noKXcdS55zWExoWU+5JwQGegLBsehkV0Z0gfEZe9v
Eq4M//jOzeaKLLu8X0t4fP21DiRVvGj7caDe15P3j+WRXdLTD0gZMTZYIQrBQDRPGPh624YM0cqJ
NLBowhtLU7mX09HASU+ScILggVqem33LLcqXGof5RMH0Wdiv+t76RkjC3Jz9ld7h3Fqp5zP+FDJz
QfXId1OuDfeZFmZ3OmuMlLIrV2QCz9XPR8N+BfeHmINf5p/SlY9YXPAG76G6nh8DdJkmX3AtdAzd
bKjAnAscAT2W92frW0nldbjcpQAWmm1jIMToI2joDFVk6C7wq2daAJx6BJxThMtWtY8Air/naCfw
uCEaMbZICoZLi7X68hfX/2QGm2zwqpj8b2G1OUtpuzYwe2NI2TWakakmu+vO+fWJqsv5Z0ZqM6cE
JvNQah6cRnot+9eFbt2+RQ6YTrHgrwmqSwURhVFZDErwMdd4XDQqfZCsoaAozWnkaRghsZBAa633
VphRCPYDprtJj53/cImTcembJcFzyHJB08J3rhXHZy7C3SaW/6UTFcllu8iJN0ZMmjKUCw6ZIliP
93Z8uzcP6gtAELtJtMaJqArHin2HaeZJA+66VtisaI5XZArb7Fa7z/YsKgNFDAhmyCKHgAClZbwu
89VBhgSy3rSqnMYFhGmy9tcH3Du2leaHYQDLHFGqqrZ34xOf6TlDFyYYXMXaln1aFYsvaK6mMI1Z
ez0W/GRgLu8nhPMrZnTcYzrye3VZMPh8aeZbKsHEKYRwwgy7dVw7J68qeg7mTYlpITpXljnh4LtQ
s7SiJZTkAzVUu7PzFniYu/Q3v6Lu1Yrj9gMIYVhLutJNQDcRgLQdl8hcIAiS1TBYShtfcbjGYlIA
jKsl+M0PVfxeKVWk8fLpcTiP0OCU6wqAffuB694Rdf0Ps0YrGoXSdWIOM4gfNuL1KBqC6VzJKXKM
NaQ+CUR+CuNcBfivSrjWxRlRrYdxD9nouBllUuOrzfJcqVXnoeVZZKiwS9qJrkrKrhslM+x/bp8O
NTy/fFCAkMzkcRmCzTRuP5h7njaEr+74pjgfvaUn/NoJCDaDKIYP/Mp5VyMm+Q23NwFPz6IiNff3
bpbE/e20/Xc+pYOOWLKpNaTYdvd1JP+cSa3/tEMrh0+fGk6WjVHOQnTg13PQK3y/EkhPWd4ZnFIF
sPtCCRZmk4oP8YMR3cIrMKIImd88qTMI8PvpRVw6xj8r6cXwe/kQVDobmtdR4lMiQZeTvkoGysZh
5HCTgspGbxEs0FdSb5ldH83EjcakXxG8GQ75ZaXbtsoduvylhfcXBOpLqHBrt48EVVt0RWpf26QH
Tg2Me58VWhYJTlQNR/xEtD9YfIwMoyYOL2LQ8IgoFkJY8yqWjaQypmbsnZ2lXvZXFZacklFbPcwo
JBWQPmQjK/MpJgxKsleQHztP4WO53++IAd3grQqn7EbY0tXyhR53lXh/wYNC2IWB8em3HHh9xTwo
oMi4CvUKvjNBe5IUjzd9OXj2e7X3FMwN7dk1KWLSD/BRmXvgX8HV80Wm+ROvcyp7PJrz4uWhqELQ
X7jvAbntxFmYCa/t6NFWJdtImTybq5qU78nIdS4p0ryH+eFudLVH35T/tlUlzU1C8i93oHJ4sNql
YOY3hiEzjAfk/wKZ/bfB+sQof0wNjuoNFvdFmVteUlzFGxwI/fPR/qxhaiEfv24NddO0kgBqr50/
eVwuu439X67jOR9bWy//kPbL70VVfQEbNIi7zcn2HLYNr7hY54itZ5QjQE5k5yUmaXkzVUAvvhzw
k7SNMHoV7KnhYtlOUmrgQX4VduIfjcGEAiFLVYjOEZ+GkK1D0OhhXg2N1JwypG9TRwq/CLN68bV5
pcqW1Cn02QTod1kXJrWPCyGKakPb4f1Pugbb9Il2WLJXQLeCR23lGP6Y3dV0suDMWDyiBaMKGXCn
8YrNnfsVaY25alRqoFf8dgd0QELvB77zzVpsJYgR2HHy6PZohLnMel5X0m4byw86OZKtUnYvlxwC
66lysO+vIGeIjoXV4c6w/ATiW+cDV/MUafzAA9bQ69n8t2wh1SpB5FY4qiOr4Kxh7Df1l86SM2Gg
kRYT2jbh0m5BlCTskVikGLGIF9QrPilXdR3/mfkzitMummV1IZgIMgCD0hWGIHSLMxxeqJqNJY//
094AdCp4ZdNc4KLEN22Q8U9wnyoyODseYUjQZThb7C6bN8g1fZNyCecsFSdJvNG6vOEA4JhxmLUC
FYddQRna6Nf9w9oMrKqUnot7mhxvdUdttgye3/sGnWyOU8AVXfS+J2D5gIn8oeag68L4K9n+62IA
am0TQha0yQVa3askAwZdVheryR36qn5kTEuiXlrZl7wBO/+2lzTAJw88R5Ih2auZsqt5oXlfM7Np
TbalKbH2TldatMYRj3/GSk/WY7Qpq9UuUfq20Ne8fjhmDjP17tNfi1dkwbW+FXXNibj83/H2kC9Q
17ZzHhsM1uuM6aDkpm6IsxNk8NO4/4P+nl4t0jJuR6bsKQ7aFZMuUJP/OIOwYRNmyK9oSpLQtOr5
0WFPWgYwQ7Bpq1F60ER++C0r566xU8veAfUX4cxyP3SbCjfC7OVqGnDTlNUgndu7Atj3hHHqHeWV
cs+hV5nw4ojK2Oj+ccQHG7zFGEioEW3a3JpUHKWf1qvqDQi3wUru6QhQoo0UoJ19vQUZL4uws64W
yLaPuU5NThGz8ADTEs4Xa/ocpDOl0yTsCSYkBxcoy0gnoOnKS42/mf0LKiVjNwqgJ3nak+v2OJIR
lvpltrdHiEKEKde++qHc0ON6S/bdsWXOD2luGIRo274TBsH2QSs32S4GINm1WadchE1dQgSBVBSY
FH2ZNkPLBodgqSOCN++4shD++Aj540Vk1lVH4c8u1lPM4hM4/g+PAN9k5rzyPoLH4l4TQHtlFQyX
dLMBKdhHxT7JOs3WjIM1U3MDp1g4Kyoy6nHZhS9b/idV2WKY5S4smJjbgN9LLjt1/2yI31VWbH5v
ekxB4iSK4O5Q7pd0FfIFLqIKUgLB5u3B5oWi90aXt9BYy9xSdHLFM/uoMfepeLR+9CQoRILQj23R
p1bjkGKsOdFWIg4IwGIYL1xBJBUd+LiuBAuHdPjpmEg3K0ukyJ8K00d33IpUiN+kkzxOKbCNNCOG
5oEFnznFp/NIG3nCHPNQdTbICYCFhYT4QsRt+CjiFrDh9jPRF0agt/A2SWAerHVXOM8+Up8tVRDB
nSfz86Ut6Uhg5dQ45xbMZWm1dER52aUxdf/7H9dg3sedf3f+305STitbu95cJU0Eennbs2+TjcQv
nAiWBpsXFlvjglIxKCvGAHGtJzXWDLXKwxYjlRKZrzmbHEqZgyywO4L4Ss56RlbO3N3XBcR4JGRs
ChxrvH+/aXHlDY0lLPIEIO5afSrQSJsHdX+sxhqhrBst21tNuPWCkR0Lb6BZvSaCE0l1KgZwHbnP
4HiM3IcbLIeM7odE/mH4obqZ7OcsJM73a+oVMhxqy+TglZgXraak2vo5Np+qIfKe5+KKp1PbadPC
dL+4yg7C+DU9VQGXyVBRxNFVCdXA6cDEgFf879nKitcf++2woKdGydvPSKoshIB+sQ872tB5EnRZ
Cf4oU/yKxP28kKbs8unBlZvxLeHGhWmhdYYeXZl/Kx05j8iG9iGKQV22Q7yreDgb68fiV/gEkvRe
zYB258ohIhEW0y7ZHSC2pNW3f5NpkuaLoCZm6xU1kUu49VeTisl0qFvsvczAcjoCBrLfCu3OS67f
KAqGE9HwPnuq4Te6W18V0LnjeHjLGHEuA993lY4fZdjM0wJQtx8U+rdhZTM9EI8glmNAMM8ZnVE2
yYUrFnhFMC9SsfJs2qmPke8cOsb9L5gwOyqjoGN4pAvwWHUlPjVwTiDOIPlavYAUAAsQJ6j36qXY
olZfyVR0XzR328qiLTLw4ugFaCypH4jD3CNSCamS4kxIM7fPb41MQ7e9HLLgpw3KMfpduymmXYms
KwTffrfoDwQE/T3+IRVS7Frs9IZXar8nqHS1Xi0YG5hDn5jQ9pK9EWahU8eqOGsqlfSPRjwMfmIt
BzW3jVQXRvJwsvjMbCjq5x8s7LqSOeKDJ4L0aU3VWWIzQQfKz3FVO8GoxROc+x1G0aP310MExt+3
NTrmzA/yCVmu7VyPfc3IMyHfykUVWn+wB0dtuw2rvcnU/QHuOkQlnWHjAsUjlL/pUdkPN1uDeV4u
2wljJTC1CXwkm/RyFVggiJEnD0yAPfBV5aJo887yiDwW0V0n8Fqt5/EfxkBL3JqXIPmKOzudT30g
KUJefL3Bdne8xNv+jjXKsAvRaelJccZLuLM+3nV65QX/wf/Zw8SRiPLcCvjnx0SxWQlfd5w7o6B9
SiDtWWvivaMTEh5Jq1sM6BRS18T2ijAyQ9NeTpBRA0K2iUjg8WAHUky4LZMFZ1BLWhfAmO0yTBm7
0NP3fxIeX07D0kh7SdsY38eCwsCGcxGYmCxMJdSFzXiCBL4GigM1WcjIac+LrXoR02Y7YWVZP9Vc
dhMqaG1BDZDn+poXI32lKFzcpgE66qnt8Sw/OhGc2jHWXHmF7EnxwSjA2qBHuZz0kiaTKh9WWlKP
Sj2MpFni/zLzFRA2nL1C2tJk8EXx+NnTGcxbwalN0ucDF6APzyo+BBEDYdsDgESUZDrF4+RqV2xz
MIZbuiXI7fmAIjE3oShT3CTNjcHRdGnyIVCPF1cOAAqi97JjBldWmgMD/bQf3zax69bSfRsKoXM0
tT+C3IjZdvAI4V66OnXOft4IeWohX9vVgFziJIj3tF7QZpYS47wUUHQPGgHHwCcEDmSh74v1PJx9
u6L3Ak6ZpFjdRhvGqCZGYd38GBk9gLONAreQ98Sv0kIQSp7LF0mqBvdJqSCnpVv4QK2fcn/hmmeD
GlDyI1U1HC9nBtfxB0OlY5po4w7bcRc9YuLeRo0bElGADgH/1Kmb9TJ1++UR1ux9mBY9xrH6xIR3
j8ZuqTkyDrGvrG4ULo+53o2TI5Dh4ojOrwRrUApq4Hn+uETuoxGMODkhpnP+AA2GfRIwPipd3aR/
1C2RZB9GiaFXWjOGerZnHBJtTtIIC/+A1/vdhkuqGRd+D9gOznCRlYGXUZQqXH7p/jBi9aa9B6ff
4cJnKD8JUq64NDELzlnkmnk6AJmIxW7gWcVa364zQ7FcUu0MHNShPhx+se7AADOQw0lT3NmVkQ8+
eBXckyg+bVNanVhvWf9Yh9tQqyH68eB/fW9V21pBurrBewHADBNiJVbAttiCNvjTzHm+26pHqiG9
XTiQ2u9MVmJFW5pkQpOQ550EaJWIYyuGlV7pHNoMYE9tV1mBOGOXuEMhArRm3oF5U0EvyyOsBTAG
a3cTRRfCHx0t1rxnixIJeb5jMBRafCES4fAawOEcJ013BAOxXMn/j/1A1UchHcVb41gcDYZ48d+k
g0+jOOe6NuCly6tPgpS7NPKFN9EjtQzQzcgqg9BLQjrUn8DFdKWo3fRClCJxEXrmyHVGNgUxJAbj
aaguW567XQZMvezYWOuHWMQ32XLouW7q6hchcb+LsmMqqTk1uFW7OvrrdXwj3fCLmH5+Fm7LONP9
yFentDnZ1RrQ4MJTrA3+0PkDt4BFEQxkl5sSn22UMNC+2WLBMFkxPDRae0+wINFbKieacVZUkgeQ
bsTYO7EJoiq9uF4MtjmBJqMT+6yspDpLMQhkmkVkIiDd3QoSV4VVGAI8JOOJM2qINmszBuPE2CpG
VQs3vIlKqV/vqMocdj01+LKWSi0YKyKWLRj63Bq2o5IWjXWrG7PBoArnpG7S7qwzIUxmmmotH73g
qx56wdKIbhFcoLR4Mnf891T7fqZIAZfz27vJH70l/EaPZBekBEqKPSb4Jqv+EnU+o7ThgJ0FjdRp
oaS686zCVWsvZChtotWLSRnAdmxtne+Q3GSyu8JQ4OGnlKbuzx55JgMjoL3Mv+gKx1aJU7zY+RkG
S6Wf58vo1/dtcoY/cZJJXDdleEXf0skCxTEadKk0cIhEPyRjfkk4TfrcmabYcdcCO5V19gildm9k
u48ho99e14A3SScgp5MYmbQd8jVeBO93ExkxCDhpx4AqCicpk/wmlaLVyCPjUTh9ukwQ0blpQhZj
u+wimuJ9Or9CiqrwzeeYpgYob0ggoKMBk3CFNRKSIhxHJwI0ApZEhhGRM8SrZ3gTwpfb332BsTh2
Jai1zeCsl59pbAMH93xdSsJ/lQd8hBgVYARLO1FSdX8nLHqZKaKPvTydNJxXmdAYlIjo/cHWgFNU
mBj6Uyu98bVArV8AI/qMj0bV79+MophJ1icQ4+KyI59gIzN8fGPYFnAvU8QTIYX7GMSM5TB/qVt8
rdqXhIkb6N1qlpiZzsjxZQQT808iPC0/vqq5P0Mmqay1FO1GJFY+05hZc+/h97U3wQFsvc3Pdji+
Jt7iNJ0thfDx0kQDAkowGBPCofWhZVYGjFCDeElpBAbPKw7AJozU37O15VC4QuiEE9yFxusZPbVX
LXc76A0c2uRnzmfDAH6qKr6igUeiczjSQLhA1r2sxtIvPyMZ/cYjsyPgVHYdXqFuGPTZP1mLT2Hp
0cF99OnuWiAPJX5N44qxefRDg71ozfm+H4uxot8Uu0P6hKMLCOcawyCDZv9Fx5ItTtWvX4q5ZfuU
p9XAU9OcBdG84X8o11sBZGeGJIUZoCdeqoRDM2+1JCSWvitGafB3Z0O3Yw73Hgs4RxKVHMQWEY12
bmKeP4rB28rSp7ebG6C6mUgHX8DKqK0wWiJU492htaY3DgOtiytbFhCeuYQDyZOAzNlZwKeULaB8
wrSo+GaPZF/bPM7rxmw2CMEAZKqtVdnr/05qQ2f8XPrT8AdHaCsspfTYPyH9Ulaj3DSnGzsikyrR
5T/gfEh4baxjRgmqNn2w36Onw4i6qmQ1M1lZZbe3pq4hmgIFRZTU993jqPluGETdb6FJiv8meFU2
xZSOLWteY7YHDxR5HR/TjCen3b+osta+ZQTx7bQDrKK9836PE6rWhC8AzepTFc/oUV4AFRph1YNb
TNiL3iWQ4PLjyEO7/FCv42azDR+fNar1orZb8xUiEfruk4wCnEYgI6Odgw5BMpG9UyIc5Mi07A3I
luPm6/FoQJt7QmvajIf6Iqh/CFT/SXB+AW4nHa8amAdPccec5g2WbH2jbuHGdwD+si2L431CaFIo
b2k8ZV7im1UxYkimf5LEa3VatwO8ZOVGPP08I2qGQo5FNWNvDnaD/umbgLz/6C/TXe4OoS2HCGHM
BYfjzo+QdJdDvPM/9IK3u7BgcIkuwJ5ZAHmV602B7IKUESUynFlqt+Yw6lV5oGOGTPDGtsOw/PcE
3jV7PZEYQHuEHjLOVjgpjJASsYstWCOaTRLOOb2jszQUCw5qNyOvfetrE6M1k7o727dj8o3zieBH
lWaz+zytqq3gZIpY6+uwK1l9fGFVbqnpfTUaz5sHS6JU3ng77bpDNMGtF2i/F6EgotbmPJ4yV74h
4jsJJK8HVEDg61A55yQ8+NGCTMsC+axZzmZSTeoINtZMx3hfhUZxaBPsxzxsQ8Ff9of7umwddRK9
gprxh9f/d1HkyFuACuPPHNJuW4KNOucQu3ggomD8ocOqX32NWV3bxwv+lHFJrpMWW5UFGlBM0EH4
kMZn7/W3WAkrPleQflZAHO0HhtiXEz3SVkUjRZNqPRgyJ44SReJxaLC+EqnRvjK+H72rwTSpBYh3
51sNltcv43SSm2OGq0SIGmwPH2Z3whAh4Sn4wa7qa+KmvoPLX4kx2J63GpplWCDhqCTEjNO11hBa
GKekRHcNCEldXyAfBL5nUgGVUUIF3cO89G6y/BBeYUjNmSWMQHhFco1dH27MT1B7o1ll3A6Hc31P
Dk/fWlbHOdVTx8CJkNuS7dDLcgCOdF6t79Z2UZP96r894AeQxKKn3lSLtfKgVKHiWa5I5xtOdU0t
DGZ+muE0kBjCP7Gp8Jlkq5CheDxyLXuCFiI2tpFlBqTZB1ttzjgQeceq3oQssloGqoSIlR2I3v0C
bg2CY861wgw9yGbXZXZKptRWslGpyRYI1qNLvyKpxjQszeo0tEpNJJsLNeO0ZBTDsf+L3LGGpVLJ
wpwz0Yq+HnQdOMx2UXVT4LDUXoqwS/ilMJaECqtK8SYwL6oVKLLTTIr2wn1qanWbOte8VFvLL0Lf
dQjSm+ILnBIxbSSfzX288i7hOz46cV7Qrd5uBfVXCJ4opGDwwnrkNbTW1JSXUH6U+oG4ZbR5h0YV
W7B3v7iIydxi7u2s7/uQWk2J2dBgJlDxhtt3cU+cvBdaL1owX68MiOUuTBpnLz6DwkmoiTXoLpbA
/KcWp9IdcJfl9tScMJH+BsDQs7ers1FXSxES/ZvyyVTVjd4Clojask0HQfiBWCuekDBkixaKfRh0
e/eCcs8WEqSIZim/BKy8V2djzxGS8fl4IwLY/iGBg7ifYYRxpHzBS77G8X64S4eoM6pY8+8Kr7e5
mYJ24PNhpcrbFpdAgnoTgh47hcy0jkG0SgUuM7h714ndaJI/BtBqJr7hlr+tpGk6TzKX4ybaEHjY
0Tyg/+2ydcKzzQjFGg2biediwmzeW/XU2Rx2y6MKfkZxBEui5Nfjxj6X/fG1/5bK3n15GEB46ySA
iSkp92yOcBXcKsB51ELE6Yn+riF7n/jrg6tazQ7EnkvvuTi4+WPydkzNa0oh8ui0KY0dNH9XfCOr
tCxexM4i5724OIu9qNi8wgjYWDiT62Cy70bOg6DXS+RaVeppG70dwxaSaa9j+nvFhOymTNBrkJKL
U8arvckSSeh5CkLHzPHPgwWaxHCrr0k7PLdq54SPkOTJVbqJOfw1+DbZ73oSJjINtO1iWZwhmIUr
+14iGLUhqwLvOwZEJBRsOqUjJZZkejYEMrDQtsy4fBO6JsMz+r1kWKq8gbTl9D7p4NuwEcYZnv5H
5P5h7zhOKY34UXyFRHyLcL+itDlzCcjyD+38M9BEgrLsHeb2PQw5ty1kWxkue5Bz+uQ4PErFaDAt
jA79017N7qfth0j53juqIZYX1F1GTHxhJuGm0pGLPdXyGaOLJleym5qsj9fSE4hocQRmaZ33t9zQ
fRRCHvlC0eJosbBPd5vTpMfEBP8ImHPweXbEJ7mmnNGbgBvLLeNwSxs1RpeAdLl0n9KJ2E2bebuu
K/B/wc4Dwmv77m1lawxOKZMFwRXOiimm8XYkqiqc2JyfkhRQMN99a7OZl60k/RlFBmygyOJHX6B2
SMV5WLpaJzZdRZhcXZd79XFGsV+QA1KTYS+QFIZqNRPhyFkWd3Jd3gIPx0ocHeZLK7BRS1k5YPtY
r3VEdYr3EPjDM25nl9V/V7aKhbduplC3QbepHDt3bq9swg75SaxINKpN04hvuZixAbvPD5c6trs6
GpBfuKiUsJacl2dx8SfNeCnpZKd0phlz026kEmAsCyWNd/++rTqLcj9NFC+l7jVzs5cKjbyq4auH
g7sB561nE1aB+OVGWQuiEqxRdkkISNBU42MtCUqDzgJwMYchoGlYDvp9L6RpwvhJpugzF7eZZ/dC
n4ROrCNUJfFEHb++7HagDDPDb1E9S/NINh3qZD7wC1jjE/y8mKBzz9y63YaqkAa1GA1S9t/Z3jbZ
rHyqODcaQ2WENO4i66gMcoxmMlJe2ikltpjd35lWwC+qlqWBcmIxwpIVeYDNrjWQVzlKV5G8E1RN
VhjNG7nAMAsg2eT940wN9kWcHOEIs1g4yGDhwNWnjMBcVw2KzmgjvA6QUb3RGmJaeoiDbB3E65/j
537GqXXrLuU5ddRrqcVpp05FjTdnW50NZf5u4CJ/OsAXictkrlyXhzSNN0zLvzmb1ERGF846uz1b
QI1n1CmpVyHo4On8J0ohr21LUtBBHxVqNsj/La9HHXHRc/g/KEWma2XhQV6jCxmsVIktRseIE/f3
5Pz86yzdUJ3h2SJS9eZijzGx0xerewzFxyTA1QJ5i4zfDUAnf4VyaieBw2HYDCYGipsN7Hgq5ZXb
q2PaObG2tRvKrBZZJ8zZM2Nbdh9vkK0jRHyx9LkqBHjT6dmf/gcCq1Ao2yYnHb6J5gkol0U7KIXJ
CqQMkHEAP6DEbhef/g08OaELNN9kRlw0n73JD41F4CPuG1qHVFBGEbdVXCK1m8B2BMffwcvJdzB6
hZClaTzKwyJTswQQ0CSE2+p5vl5wIyic8r2EBxNHUWZq2La76Bwo2mY/KmYqhLi3jSsXyFqe1G8f
5VVf8vbNCwuBstEOk/fPJFIRz7yc6FTlngrr1exaMJ0aNxpdZEkhbEmF3JVWe3zPYdW4vMHgTmnA
TCVpM+MewxvL8kFnAhWt3RyX161wDqF77TnJHDE92HWTDPtxudCw2qh7AMpqao1RhVSP850ZVGoe
Y1fhEDIes+G1JuVuPnz/yk5OhmRH6Un1f9fwxuw099oiMoBchmqbERnadNcA6GGdiLzQrJbWRDQ6
gVm3iWgetVU3tzTgqdUDtBB54nZzheXYKCpAls+1HqA11jAgdOUZArUMlQ40S4IbmG5JGKVCjZj9
wPYoRQOY9ZVa7qTbh0vI+6N8tDsaUWQdQJhnp5u/oppSuXMJaLJdhudZE2qBK6H2LV6fbA4nIXW4
qbLmQr+CF8S/ep9TUNSx0NCPb9IEf9ySrBX0vNPi7N3Evwupb19XfmNyvAPENqXBeahHOS5Xi/6K
vrt/GyOG9JTZNxC9WeYJZdPdVV/yzR/2uIHFGz0B322iAeFkxL/uwZwrebA++y5EpqP9t9GjV6eF
Q40ved4dwWAj1+WbCeCcw3+oLG7V1UaShldD05LR904ukqsvXncoPLVrjoSNvxApCwDR7ILVGVVv
YYQeYpIfZsZbguC+t779Vn+JHbFdd0Y8WTZNkaHm+XWxhlraRFyYig6Bg0PYkuIVpQnmQgC7tpM3
H97Pph+Mn6yiTeehh4mcnxabIuSEQ7mu6Q2RMWlOpC6RAVSYeb/w+HjA7NZhtlMWaRcBV1iqQb6u
Uftp1TcqIOU/WdUqk9/F8BKGHHJJlIIM6Hp54egkVDZ7umm/bqu9LCKR6xOgmRC7iH842C6vgCUj
l/fTD0X44SsYsN+CJlchm3D7z9EkoBJp3nQRwk6jEFrbEGoiJbn5HIQy/xajJnLV2CYjD3IuSqmq
ELFLcjqdTouY+M9qotFuUymtGIFQ3NZqU+n9qmYQpKQJXjosN8SsTDVyXm5zDkx6UlFvIgVEYVi2
5qwtDZ0F4k3ZenitVKXnmu4KF0P4EZ4iIYluCpmp4LckTd1pE2eVLG/fQBsENG0Lk7WMd8HJm+of
n/eMR4JXpl+SUbsEk1hUaNg/FBVzTcmW2a/8ubApxwQAOai5g55hLrZuI5ICm4B+q81U2HdmOkpX
nEQBuNdpd0RPOC29BWWkvU05KlOaNdhR+3e7WWHjdBECmGv8k0KEXK3xFhDHOvxRXxzKGkzmRbkN
ub3fN2MEBwRvyAFXMvavzavSa1MHnIZSTjjRy93WM4jZvO+tuDt3Nhpz84J9syESnj/+7qK6fCdH
2SLxuXT/S/a1mj3GgeyAGrBFJLcbIC2HgCmnLWVM0LUesdFMyxBfNkK4b84gL8Bc8Cz+M+Xiejbd
L82ToL0607hBjKmsIBKxZT1LhtUvjgP3dROKYetzyDsImQUW0tyEuL6cS6WnNc6b2wKfd490Hjte
ESlsA+i52jQXxrrHHbje21Xb1Msh2J4LNpQTNkQGSkymtYuJH2lWQIwd7TscZIpDBZBWgvE9igDV
dddDrRs+ZMs7f927PueS0kKhY3xiS5jeGkxTRJUpdaATOBH14sXNJWeJgx5zALhhjxYls5gDxXkx
pXNdBD+FfLR5rA0CMiM5WaDF+jHFB7O0UjEdHZii9N/3IL0s4cPHofK/8hcvlJnE8Nct35k6wazO
KgiQ3/1+sL3mFkYIIWgnU9Ts8tVlCD6m0J53vXjA1WgqCnzeJOtJ1FjABaRWboiG79g24FzTWGUk
bakEn6JxAzeIxqRuwlThObYsQ/4clRxj8KA7WUlAe/F5hmK4kGXR+KaRmXUFlQfgeGNMlqI3cT7a
HFHxzPqsvPXI0sCk+5Gy0TE/1dNAQ8UqWRVUTNch8a9ddLjrk/krOdp+XrTZ93j53AiHYXU98yRp
ghTx+49WrNLZS6sHsF22EbxWgrN5+tRfN43+SHInh8YGUIx3yce1a2e7JdnUlU+R8wsUMANOvDlU
kn2T2cBkA4Jnl61izrrcZYPG4WumHuxLV7RhaXwmUSGNQ6QDBQJNGNzHvHxT7LUzkc/5URYPcfFN
VG+yxXdk3nCDQIDLirdJtMbozFK2XFWRaweHtrfLpFkuuNgAqPgjLPkSrEJTZMcAm6PSpN9lExiT
xRm7CQ6QyJ48Pj3rMs44R9SHUfg8Q5wjvUcVVdHGAhDAix097MnZFDf6iYLQIihmdCf4+f/ke3cu
PsWZdfqhe5wpOom0FsQ30EpXUR4MByqJOnMYYYKbDR+0fZipQA4O/C8N2rWFNoZHNDUYewbWIKzZ
P+9wH7RX2M0l7LqEscEGoB/BTQYPSZKxmBh07zemEuI+3011CrPbtH6sef9zr99WopA00HiNKuGn
+/VBtqWeCLCBb1nwuqXZPxbWH749um5HhXYMi+Y3ksEqM1U+HhbIQGjhn3O/z6EDdnL4JUkIEEyY
pUA3l0/MdqCKcog41ZrFW0UzwiR2M0oX46Mg4Rr8Jg6m9azA3PsI4PnJoiorfW+h42LrDU46BVho
DRTjiZwTYTU80cXz5WjWaY4MtIigmbmKBZyjaoYBMXJjVX7M8gRxrqQN4Wmvx8xPCF0+MU3OYpq/
z2D0h/VzjLMp7aeJtumR5wq6+loUjBEfNmpKON502UDUBpXosucLgYJgQ9H+WLEkyXoBbX+kuW/y
UeypZkgJpqegckN2CiN0BnDQHpTghovaniopcmAw8NsTjot8CtSG1jdgDN8NFSrRiu/wWaG9vgVx
SA1ky6VQNaosOrAyB93PNs5VmMe3zw6vAtkM1qPBmdhqITnyVy1+Hvkk5FUzgkoBP9XUOqWp2L9a
BPQAo/7tgwHxx876dvzU3MOj3B8mHlCnbGOmKv9WNpUAjRVcZpFqDdqyS4TKF0chVPTPqHbRuCHt
wvXi3VQ/LKV+Xm38fWfd70fs62k13aLVYGhF1an5NsDAHGAINQm1PLu4rGLTJzCUTaJQkuKWDgat
z25LuVgyG7pR3Me5XLX8v+Jy6tajY8t/VvB0NGA8+cUHsaosRh87pgBmd7aa8jfBei0POg24aSXo
MjDgY8xN+pLX8D2vyKPfHwGm1PGi5e62Uko4/rxUsWpbvdYocPZSoxJo78CWTeMl/RG5nfdlKAlp
EAHgcBTxMaqWuvcq9iOgP+om7Tg6AwdZcnufZbgNFQRGeMv0qGo6CI0sqIRgr1d9yLW1OohyAAKT
e9iiVoskGC9wncWSQBZUgogZpOzRERDN1BwXZMM/WUX0027ESemMKv0OfeIEcYg/LoLFyfnj027r
EYhONZXE4XIR2tIa/FY0VML26QeYggWej77XKVzvEBPAZgpOUkL+/XnLUJhJ1NJqCeliQZaYi9WL
SJrZg8bxntZLVJd9+F25cYGtjyNIKT89D3EU+KZJoFyP4yLa7ILXle1Krkhe1RKI/nxtovCTBCSe
/EB0lHYyguQ7cYGKDisQbV2GLTH0yCOdR1DFjZP4fxcRpBSI9vnqKhRsGDJZgioMWm3TulgrGG4P
LyHvNhdS8A8OJwpLyWyuAYCGk8QmoHTG77ZU18W8SBqlOqOEvNqXEFohuENbWpVLNUf33Mcuqrd8
DP71k4ikEp1hwBj1K5ZY9P0RZj6+akc9AXtTwkDrfrw1obCQ2ziydA1mbbqtSYBYa+Z+4k5D/BjT
LrzGesxzf6wMqG+V6ITUHIeSUtoAQQww3k0NNTfAg2fel8s6voMR74mwZn8N7d8x4Mi46E/AzwsR
TMWYkNeyGl6gWYw60URz4EhkIVlef/PocGQu8T0OIDvurB+wCOx6LsjHU+ui0pGZce2iTPs2kO20
S4ao+S0UiMDIkEqSgC6U+mF1hDCkHfCJB7M10exGmF4EV00ibgR4V8vCe8Eg6CwpVZZSyI/spl/d
8JkVio/uZ0vKIv0Lxn8v3P+fcWKHenyXKrt7eb/APn/n0J98ZaQE0tN/NkKm0wpSGrkQ8m7Bb8zZ
Z0yK3YxMsjYzNOHtnyRM0LtwsAC8nIORQG6kiVslsX9P5zGlC6EcvXm26Q483aZZ5eUY1eem+KiN
biDZ8WhVwW+FRqalJQtwjAdGlhq3Scl/G9it1pJpHKuXgZw51jVaY2gPzxM4qrdz4n5LpQ/+npZV
mq39KasmhASA6id4s2AhVxL4E9sVm87CDAKBBukvhhPV1FJnhMMNEKSF0g8X6TFE2fUHGPiOAQPl
QgsI8sFXFS8fF5Z75QYVzYpGW9Cbyvc6MPgCsCtq1OEAUP/z7DirWTcofbRLPOrwf/d+oEuPl/zI
Y/vRZyRBSnoW5gbynVz5GllFOpxoy8IJzDqw5GLyMNFjtuqn1FqcvA84JCclluPL6wiFc/o23T0H
gS3dKoEdwj29/rtgmG/KgxrzGyENQc5VYpPs+thHhWumiJ5cskR6pZynOn7+ElJK+ySRFaGEA1xB
Jwjuu/1oXKegCtBVqt5Gn88hZPG/YomYjGKMxjxk73NpRONlE9oh2iygPX4UOZ5o8ZEPFdGDuP0g
bU4rnkAZ2Ym8TkaOSnxN3iKtN8KTCWnAXrOzeLjTV/bC5QcQL2jcF8YErSfBYTtAAE8On7/FtFug
S4f9EfzjN+PWi1JVyFSpMgNIH6C5BgQEYY2a5XbdGsNuU03HaPgu+8FJSOuhmQWea1ufsVTiyfzX
SCAsCNf8qztTwElq2P9RYNvW7zIG4aO/FWwqEHDaIzTBOlOETliS1ecMAlf8ZWnqBZG17OjN8rwj
vShyFaPdQms1o2+6uaTldqHfjgMb/AstsvqAzh68tEvHNTxpkrZ+yUwsUZ+qX7r/SWmSzWoREEw6
LFRfz1b/FHr7QmE3b9D12DGSUIxSj2JEuj3Sp50whhk/PJhdv6HueYk1194kDAZa2kV/DBNJBrpA
XxFBpIn1KoTqdfo7SWiul5R04xna6pG0QunkYHONSgc7Wl7omKTKbo+Cfx+9dFj1vuJLOjA0rMVU
YUXJIFL5CfIWRyjaYlcX8UjWS1LFxMQJ242lhJ8D6METcdHor8uGtQp2VmmbH4yl87dyjV7Zo1Om
iUQ9ri39jykCGNop3Itr/Bkv9iwgukPtlHzJWzDNPYUvG9EKPWBWR04IBDc0DrCMZ7FviGyUiFtU
+mSYVp7EJQWib/LBNPWbBEA4qjX/O7K3nSDXEQ8R8VgZ8UMdDik1/11IMsHYf9eph3fXw46OL0ir
UvO6B7Vu9cXh0lqK2nnlFzGmx3uBnuq8MmRJowraqH/G7YnPn+Rgb+QBFYtksf5AKkvk5zOnOlHg
7/l6liwJJk0ZVvF0uwYFuMGXw+2gd9q90afNxfiFzeHNfbGVMA/Q0ECsRJ9SX56RZEGrD7u0sagP
7GmznvVlOUcNAd1LZ1PWj/KD1hB+MckwtSBinmdyXpqrYVJrMsDHZex10JlhsJxcjRRvdQ7TGFtT
RRgsIQdiloXoVoPZTKRRjdWRnRmNe21hUFw/VrmNG83EA7zqmeSKzteSm/uL4O5rjyPeNyxyUJij
4lyU8ir2dLjWrumW3PCZisi575poKC8cTSCkkp5KSms4imQdCxNl2B2Hyt8H3lNgOEH9tg4Vqq9c
GQaCDFTCWX+AUaqvDFfMJD1eigiTwdAa/hJqtxTVjtFmgmNHWvUGr62N5uaQVWz8Kjz2b8Ws3HTZ
drXi1kka9gaiWBdqAJMfPLBDBkOC3it8niv7CSnRUDsUmVAgOzayxEeRXH1IPSy+zDsXM6ZTpZx+
BxMxpGTYdLPheAJenKM3ZskTYwHV2ZIG3yAnJPGN64nurZPBnujU0EgSxTFjx1rb3tzmkVnHD2hY
sxEnxpxS3iVOdUiEE3Zal2XaPGn2LVEYAGtBVVhlczjdJ1LfcqmX5nv885ky1EOZGWCqWQkwsP1u
lysxeyrf47yIYo/kV+YZdzla/2IN8KzMQYRzlizzJs7esry0U3FCMcT7TajI8Wmiqqd3g3y5dPxX
wLB1j/xtkQG5rvom+ORR9wDy0jEH0B8B15HxmdoKGRnJ2I74lGTUbywxx28iImw0tob2uSeNMrg4
7skAld2ACtf6WQk6SOAnm2SjcvX1F+3ca7BJ0wmum1uwK5rFofHpSc/ljwntTId+CUjVk5y77Ay5
u+XkJmBptbZpS72MVJO3nTzK1G03dX1vhIDoSBIs9iebw1cMNUpKfPAhQzZzSaqGT6Gh+urLxF+T
rHah40+9fAXBjBe+fjqsCBssaxme3fLXGeTLAiqYWzLJa8lRKte1bRnYs9dLp89d7/9x3uJU10FL
hDamBHxlTSpl+fWGsxXTOAISqsnwtbpAdNdv8C0xLfd2GirssvAR3/ifLKkV6X5E/Z8NsFB84i2d
Nsce2zin967VV6YBUDuFCRHrbEKO/Uz3EuDabJxh2freXTiS8eXqRA6A2qNmcxJlwBLQnGKC2gFP
i4BC7J1W0djw3ZBMrCQ5KCZmCTrPbSLRAqHQ902L1NzFlSDLd91NYvQ/5Hqo2ifHggf2HtWFgLpw
RppWP1op8oVT51zSLK3l2zLBaADZv1ApDbVvp67kKB1/AP+87ubHx90rVugzf83YTN07qOMymnc7
3mqxWiFU5i2HI3bLpxU1WGV9rBwOGKyTrFcmmaYO+2fceQvcz5GthZm4UAZukAgC6fOk2YqXQJe+
bJ18xvvsks3qZgjMaz01VzZaW08yd2N8nN6pDhKCj59n9dvd37dRcoaaJ+oxE7sfxGeQ9InfCJcF
e8wnw6TQHcNyXiENDD/Plf4Pw6O+G6vwtdfTt5hBYCfPUhqAswmIo+pbEmI9VrqPsN3dnkfE+08h
YeEgKXOEPMPEDSbPy35NFsE76zmK2v1uSE731wPy/0QbHJJ8Uex/x4D+MUetGpcbWIg0Vp6naQw6
ql5J8LGnJNLqIO8+6HKGO1dIc2YTFo+PrD0GwMkNg1I1DOqZqaAdcz8Z9mi0sT5TFjnqTS/REsU4
cKrLjpvvEkLmGuy6nzyAE02qtS3S22Z/aPASrxJcdJ8VSa+heoZ9HWg8DPfWKnnRIf4gkhyYuhtE
sI7aNXOvlepd1+WIrQ57kaz//xDHDVkzZYCCstqHbCwLu8jNtFlbGSrzEtxDWaC+A3T1RK4Op/Xx
UO254dmCoxxwCozuSXIAe1JggvN0YEhJn52CqoJnPFE3+1X34+jIUjYnIHH+j00TGNsSxScdWfL8
SpJotj9uJpmk8coUMos4YniT19ZWB+1WIZeEVGSTQd21MqFsVa+pjNf6z22M0Clfsr/Ex4IsKzGB
T5Vsvwte+RHWbLn04gOH7f9zr3DR1S7wzehtwPZLS4m74wBxYiPy5opmzuMSSJLK3+YAPXt5nGmt
eZ320YWdVAxZFl3Nx73bQInvG/qZAEo8CsDjXOlIXayHPPabwCvQ+0T+Fj7L5xQEctzSyXGRNZAl
YDGNv91doaPKLrOo1wLtCDEvB4Bg7g9YEUrxYKIO3dmwI8cin7O+Wfl4iC3PmPgKtO+4Hk/kqyWN
8aPxMHjDumdX24Sic6G/7odWRlxGL/FqrcExd5q9O+s2LUS7/2G+J29ZvEu+b/YKV//EqU712j6z
ruaR+kcLwTQxgeSA6HJOWZl3GhLfSn17p9qjlmhvy3rekDmcFvXP8iBlv8tSnrQXlQGMNQhiHLY0
T3mxSSWmJWDnguqUYZjsGkgVmrltoeb/2x93EEUwnaQevEZ7PC9dQ41lYk1B2Z7dz0kE33h2QpoZ
imncuVKyG/TGIiTJy7HdMzdny8/s/dJObtT3rxWoAmDIks3OKFMmPCxjQNSOxuMMXR04vva1UGLk
ihs/M2DMgxnR/AhWVUWUpLq20sSCsw9NunKhsGo2gqYvPVBPnxjpyjsjmHbtmHqQpEhkqtZZcjfh
uWjSb3aD3eAAa/QMlICKvtQnGyz4z+7WPCUMSAc93eYiPRv2C+aIa3vLr7jMQYz0LJCgQOe3ZQQj
04O7wpqmwAWcPhX2WnW5629Wc6KVKS3XrTCVUx8nvlt8UAPbDJEATsm+89ghrLbCVFeFZnOo4D1G
IhptKcSzfBJVsP7oLALYHse18Vrvn17lQl9+iZ/x57xyPFngqptt7HC9T3OXdtEYEG86p8OHQbuX
BYUA3KZoVeW1rtUCSW+zFvx1sbrcEpPV2cLzzxZzoyJb9UqzeOC9DlpNCb/MbeR5pVROy4/hD5WI
mzd60y+vgwxNviAuCSEXS34PvLt+RCKpYRzwavHaTDHkG6o+NKCxm36gc36r9aupx1+NFlPyRAOM
NNU6QZE0ZXWncEVaFmJgK3ua+ocoe+L/ooghkk7mxxCldm1azFH/4de+uDEqFAle7e8oFSF274VB
MBuC6H/5giavkJVoaKYUvgGfVQtqNDARaDa2+s6af1YpHSn8/chLdZ8KL8aXNr3CqHdKPu95pDBO
ZlQ+ym/nPdeeolV1ZFrUriLwb16wq/a8Il85dKLR8mDSJ/9exAMz2gIUoHtrAQadSHu26zeu05v/
7OYR3yiTvPMbZr/9IsOSS97sOPtQ/JxiEI5WfHITWSpGkLqh+WlxF0An4h22xJnVpvb0QLOhDiLG
UuqMvGaLqKh+/Y2hSjV/t4FWRlI6W5allWb4gEqR3Mo6vnB70azSVu4ZqerrSiny0lwWiYuWnen4
/JB6putgb8RQKHpjNvZklgK8XIt5/rAyYsqUWxu5MR6WNIkomEC0oYozXKZfcX68yi2Neyt7z3op
K3pZ4ix0CRjUSvCEf6p0wc5JNa2b7+eXvtE3YR0S+t+BDSccBCR+myM+4jjHozH4dRdtFJMInWeT
gVWtGlEnAFU9wInt3dqGoycU+oiW1kuMRDxDbfbEw17c9pzqnd28ER933CM8KQR6qCQ6CDaY2K3d
zRr1QDRWwhYXWA5FZQK0kdF8DiGwbp4AUMuMSrmk1tEP8LZ99+XW1T2To4Zr2M6Bfvq7PN912dcn
18kT3dyCJnNr2mYX1WHzkRyLhlSMY3dLblNX9FuVIYwVFjINMPlQA9DVWqD5mt2MNCLH1XKBe9db
rxpg93hmkVGkSfJVRJ3RJ857hgkn06Tya0Nk78MajVpjfIRadwnJpcc+fMBZo6iYwk24xqXmDdfp
OEwamL7tMfsqKpAAh358iI8RjJNwR332dSkGM5U06wyzbzv3qndML6dsIF4h8e8HDLrevRftzIWO
AsUZcGNwBP/XSNBH5MZIaWm9oQXhc1VzOeiTXJ/Oi2WIF9wwB55BMh1qgnfMslXh2slkGFWTo7Ip
Jd+s1asyydrzuInJLDFVEFV9aSIPLU6z18WKWYiapN/ee0lZxM3O919S/n69nEmcglissylY1Jiu
/08h6D28OkusO9uskH2G4E9ezhPtDYLBHQD0sxxT/rDlpe9PeLKPFURiLUDHnBoMEHoG5/kB/fXb
QiyitfFfv9AxutJbJ+/nYzZ0l8gCoEF0rII363GTjryuoxefuTKIbgCS0Bye/CH6nOfOViywSEwG
LiVNJZH5dM5lyX9yH5FytyD8mdf0qy8iQ78vVdSXFBrQ8y4B0obiGw5ASEFIFxvlVRo2mMlr0i6h
Nj4Zz4JwzafMReTKWqxrIQv/G6obOorF+Xe0QEGDaGtRY0rW8DPVl+q1VIAfp/lEW7wPMM2VzUi9
U17OA64abpCPloXYZO5lXX3Iw8MPTA6lb5MeyICRb7a9C3lFf5a+pljL7bJyDa6sGZM4CqUR21CX
6P+sxP5gqC/dUHZpbwDS8VlO+spL0XRIIxbKv1E55FdZ2OIKrqeiwxPyFD0aiWw7oyPZH2FHaoJi
LpRLGI15aa+0OJcOVY1OWKTGlddYV1E5D+RMDasNNkG+GOV4I1wwylWaD66y2NL6UPDrFH94EPcC
Ff8RvRrwpHLTIt5pw9hHjD66gY46KRA6TDfOTJ83wz9wNZSWCY5Zi9CRf6Gu9TGb0mR/qI404lhq
l/e0nYOoOApemWnHjKRgJ7PxFHxayEMlYQD5Y2wPeotubI0uEPfOmGTjH9J37ky5jdlCn5Om2qxk
/e/uqeFp9DXF4Sbo1JsPSmE7s6AF8yb929GhqQa155q9utBWGhiAnYJBBJwj9VT0pdsbtyqQOACM
B+KHGOUTGn5SmiYXYwNAwqyM7yDJUcU4xlJ+4NbgX1bQkYaO8PvH4ZI/rHMCRYCd2Oob+A/8wstD
QCXO8wULedofu2Aojyn/FJJgM5liRfd7p2q953AmYvuzDBhSYOr8B3eJf4URtg/+AvIUhBruBwac
9cPSauMsdrUFd3hnQNUh8vUqzhcqkwaTF3ZlrNHM/w6Q0Vl8pVGXMj4kgHJgJWlhuA5MyxbA9YgP
a+jNHv4FOxkddQc3+bCmpErXr20J4r0oa/pz/YJATcaGM1HCU2VQyfC0hQC/7plcNjZ2ZGJbu5DT
h9kiXqOujCbUVZhzOOd3scDeMbDXl52x5R7IQeLpKAwL1ezRf4nidVpoOgA4UOdkciUyPO53B8UO
T6AV2mTLVsyD4CnYoAAcsWKKGIA9kbsHvCTX4gfQnIia1ZSn7UYQoJtWMXyQOqR347rJqueM7FXX
BhRXZZgM0WH9GREt4AbpKxWj82iZFjiui8slocwApOeJdPgVB7ar+qfGT1k80+01Rgb2Gzz9xDSP
cikLEYu39zM9MbZ03Nf5pwMtDq9S5ZUlsjUAf9MurXouJC0evVSlsejVjHIIvg4QYi0nAl14FVpV
6IfdTazRDFZsRlALwLoi7+PbOHQkqXps7bGdA/sZZCfl6E50OrVqsCNlAnILSyd/Sq7BXzfAI+ra
bZ/JBLoQ0iarjRbI2i07Vl8uohn+mCgWS0+URZGp2398bi44alPvIGSmNXkjBnM8oH2y/4Bw6xW3
13ovuB0C/Dcm5UkIMErS5Sk/gsf0elaM61qnjwFCPpD76FVrt2vx0HvS52SSlSwHqSzvuxDC9WsQ
EVyYEkumf75tbAbuMwqqF/Pdj/naZ1QIudGKKBzfiHe8yqW44KgCGqxPdFd2gHpggmT0a4vOWhp3
UrBsinrvmnFcZlF0hFXthGyB6tBBoHhQWLqhdonLa51/E++P/lNAoQWBsK3xsV+yZyGJ7aDamw3w
aRsdJXjnfPE+HHxNztnTAuhtxYU0pHZ66uZo29yjm8Fp76vqe0s/g81UAgpvqNRwpKXw6mfFg2un
q6OPHccA3PZI1BzfVwYnnBH6QSZBwOGL0HqbB6EPvJnPqPYaxZgs9BrOmfff+ZvN/j/wJzMxlWED
XVXPwEWduS8fOQcQG9hj4rdt7bdaWxxQmB7SAsp5Wk7H8o/sUb4Xg7SJDIU/zW+paQ4kd3nNhSpv
ruZej9Po4hxi9cGSEEvWREADpknS4oYf4t6xY15/OnDsJrp4vnOT1oNXiNfV9Q0lOEyoMPgtMSuX
je6VLfnqA3c2tSKEl2lYHptFz3+AFHIjINx+yidXv37KntvbRQZqcSHZd/J+0M5hbzVcpH2AUYum
EcP5HUOtSCLki79he314BQmBU5icZKJWk0kScJESMcnI+XIWRdmIhv6cJhYr//bTGQEBmGJ3nC0t
skvnV2DbZMTr3AeWw20aRlh7WLbJrE9uFti3QB11q+lNFMMVTVfQNHt+u6DDq2bHtxEvPWukqesH
ZiQamzLA+in6ZVxQSeW3hHPpbuK/RNuYv9joFwpyaNiDUEJJVpy9sOb4ZUrT9h8oQBsHlQBJycuR
KcUnKNUT/pckzLaTwcIeEknUBDztItnpOHzfUDmTEwMbEQOanf6rYlCeWMhZZWVOGzlcqpXXtXNV
7el49q4GX/gIdmqQ4ZABSWsbMM5NIl3WxU3O9lRXO3hAfsaouKX7n+gj7kLzK1CyHIWxHm977MHC
3CHIuC4oQ1Q5iSqTga4A3xbAisHnT3Jc6nn3gghVWD207UnsUJtosbwKyMmcCYkOYOpj9IhCnhjC
sIhcCSWbd6q9LByqmDFLBD0B2D1dsCC0ichHmXe8IHveeSwnGlJfQQF1Q5QJP6cepC5NP1VQRDVr
zrt5oOeyicR8e+kpMVr8o0S/waxoR4KOKAywWRFVoiGKyGABR3acQ1CcoGcI3ab7Nk0/x8eILRss
IAkB7HouWhzkhrNbmL3EeDtrI0Chr1bd9z6ZVjuh6QRKUwTL+iYvKsw2Is+J9dtiNWT/7gSFTeWm
KWBi8GbFOgP9faAmoharMd1xWN5NSZXnELYBPeRp70sgkv19P/RM1kIHsF64p0+gYh9Xbul17Uim
T0bMc3MX2xS3YoJsRWERKf/l6L/U0sfHHxR/T6t/mx1K4WNelsDwWRAw2Z3s98jB6QpSDDA3OQpr
o/Cuk2nrhtNhed6KaK9TMkioH+/YQZYyvrmaBQ6mwPRkqzcFFpNywffsbcEiyMAawyvpvX84EVpf
k0SHHaAkXQJJVnjvzBtBmNI7YUX4ry4/zu4Zovf6oV61QrnJS4eRqsZKI4wZMT91o0lNIdnd1oqV
bCzKkZOVKt0R0ta9QBSXw152RAAS62youV7SRnZMg0ikLlNi/D1SW4Ep8FXVyZorVG0y+f5rMXLa
h8UWmEw47NlEKafK6GYtBauzGC7obDJogHUJV0KHhchbmIEkKyZ251kFxuQ7u+A0nfbodfrJ6DrU
S2zR33VlsQLPnG4cVJewBkSk7RiqobQmOBwowijCGQyzsIcNF7FN0Z6l9A0gcLJwVUF2k23gxyFp
1Hs1ntl0Z6sDbobNDri+ximCnClhDlVFyvk3CflY/pQsugoTULAtn7n9jbKx3hcSVilzQhxEnaHh
CK65e8ld1kMubPidmNwoEusJMmjjWhiDOup0fqFpAXvgGdF6v4Cry8Cg6BRxI5TD8GXLR2lH/Sup
u+7qNlQCEtA609bpTplKWSLP3tK6PJlOU94KiukV9LegK25iPC+lBezs2+xNd+ulrZiDJvbcYjHL
zNKa/ofYERPjOexNg18s12S/p0z5rKYSai5iDDaRtby0o9UAzYFRXM3kQyAiyyYRjB/CqMVpk+9I
S83loEtHCLPwPEzIMjBFePiLAUCRvRVCt/bo6SPLnrVMSoiwiDvUwE6CtKWT4LfYjTX3ASv17Jqy
Rj+kugjXB6UVlhYYIJtIbtufJNVX+51FkJXTGfCcIJxZtKScLwuhpWu3Uin3PZ8ptbR7Dvc9upyS
OmKPg166RUMWo43SBBhooh1s1QXPjWTpeICp50f4YlWaXKm+RW+GIaISPgxHLZU1vM1ICG5AlAkd
2cwl5lSkMA0lsnE+f9GkrU97M6T3MHZd4e0iwNTHJAeslK/XMRRZmvwrOix+XfR/oFMuHWmICc3X
6khzLLqNHmQevNPNmst3NmKlPyf/EPzuHZ7ase7bjd/JxfbgmPdgN8rmG1kLyk19P5OMowK8pyIw
8gFoLdYw4aQpYPT7LANCFkwQ9UimsDDT2jMlHWhBTRZerkY2feA51jV2Y/xfBPbHYq+Cw+5uC6BS
Jg8kY35iMOamcboq9/pWpf5DutDCSJ6CQKEV/aucSGvumSzjo8GK2oG592wVxpxdSZ2ouv0PylxD
VqCVagnwbqnzEFObBHm9qqIbxdhzsfDTcVHmjvdVd4ts8Uvvit2cOy12cLBOnEXNfEOzP2nu1Pqb
2NDxZQ0HEYSTU4ilRZYCXDjwdysmOxiSJOr2hASZfAyhuaMyuWS6jh7e2cM7Vc0Pc4nI80aGx1Vh
t2MqTKflb0cEdODEB+m0yR1LvinYJYMx0quY0BOxiYecKnYd/SMDjMx7sVPfEDO57+ul9hTC2XNw
4wwlRNIx/GY/b2Jrfyv+lKdmIkjgenpswMLv/zCN6B2k2JhlFcLmqDlB1YzOmf0PNFPc3G4bAmOT
Y9Y0fU7rVvEI2/QR5DABhc8clrXvlMCRr9Eo6yKLqBe6lk352jutDUcMGXdnLkcIJJse28fBvU/O
KK0gUHoh7YfkCzEXLFuV+T4liA+1xHBWjKfe35nyg6HxSU/Rir742rjsZ9i1XOeIZKpnWBw63dqu
rEIOCWrcb9uDPQjiOa025NxcY7R7Yf/hKpkhKc036yzdotwjrIab3+7agQ5oGquuDNJSHE5P+W2q
PjoflfqY46YSvzXGb5+KRCJ9PByobHBQv9IZUV+HGGVWB8TBjXM2M/RPjssEQTi//vPb4nWAjoEY
riq9WuDCaWaEZ5UQlGiKJSrWZHnZcTrtnGHpsTyi8dP5XFTOBVsImwXlxBt7mzZ3NViTUABV8bw0
RttW+PAbWGYrn46AHnZajyZGy0A/nwiBivhAH3sDta0p7lAJX40yELMNPJDQcKqgfK7hWcSfoCpG
Wl+1f7/lAU26g/IBjhGaHqHRaUfSOD0XgIcpM7z2kpP1O13DfjLUCHzqIMc6ODKJJMEC98cIh9x9
M1f/quVKvzdbYEUFbcyFMKgGppEILJyuJuQhJEF/cWgsHnxNW86OV7941GpPTtbIR5Ou9VJn6d5u
jOpXYo8TXqBkLBpUFwJOfprHkNtGuM95WC4x2YYYRCykCQjgAQluBIRf8mX8bXKwUNVfN+7EGcMi
520P1ubQQPS8ZW2BnHskdaIk6NSRpiHXe61G5W1K4rRKGiTSVSkQ9lQMXHeHgsuK/7Ogym4wfeyB
Pa6zEpYrhto3ONfuWiGvD9yKXYcQ3C/1CBq/2+QoJBJyzXKBcnp5vBWCwYrdQZFIZkjN8iLDTQo+
IBKusOSV7l9HED9LI8xpLKvKpBxG0SFPnv6VVJtDrm2nP8xjgtk8Dx64nNus9ZLEgScizJ+gELqZ
y/41kmratNXIj3jOe2O7DS8xgA6IvtqsOPeuQKtA8S2JSQv/Hl3hkLY+fu3FE5W+XGHZBRCTrsq1
YJXe7kZqDOKCl5k+45e3+3Wa9+cBdUFEedbfX1OybsKB9YPbWXcnq6DjSc5m+BdOpyi523fEq+OH
SYBObWukAK/PiSyUh7OnItemcgtyrwYu0TvKU9CkICuM2f6lADZ4EwrhYtV/9AkiQyvJsGAzRxwS
9/sAw1OdMg8Jdrky7eLxnrVkIeTDPU3CqGFKl7NPP1x+yxZJ3M9tJDh87C1FvTPxQ4PqYh/+E+5j
BDZJkhemptBdpUMvuhBDOyWmtAbKx7/0GbdSrmGG8MKytammB7L5r8VYmpBa7nPHTBjgQg5HCanc
KJsrMCKdSwKgcS4lCrVNbmrANb3lqgiMHaXc8pLgBCSBcVIdGJGWPh4fBFrwmcbuBJ/TQAk+8oG5
ntPspnqcmMA01tBM1js9UmrIhH9I5/9+CMF0ZmfKQnNuBYstdPjw29FVcfwpi+WkLCEhLAcdUxId
58Y3AWSz7MCQUonJRZrW6Bm1rLzmoozupPID3zdfOh9yHY/86WXMqq2mLFHuWV4YNWyh8eF6LL2k
XPVtQ1fx9EMpKBgq1wUu9tyER9Kl97GrymhDxSiPPBPeRdWNExj9TQhbY61BpfqAOh1IgKGkXAPo
iuoWymW8eRBNwj/Mzws0LHGmz2U6rcpixwSVFmDS8M4d15kzFDlwGkvVM76ZZN8hDJJ+fmX3srY7
DyzMxXcv7QLHoBcs02LY2vSIJrWR5iEqG+pEDL2J6t+rWNJv6K3up6NNHfcvDbkhpvSxD8Boxz4F
iDOMspZIgruQk0jTaFGsdty5DdGpJqMdVaysLl7RSIwUkxGk+8cXlR07s64AgY4ku6YRHP+NDry9
GO1kIyvnE3x/sReiCs+b0kUzpx8fhz3a4T155ylfhaeyPhx8d2vIXRaI7SYConfmcA6/8kKRyW0l
Y3HF2WQQoy6DAcNjErTM7MIg3U3pYrCTc7IWdvh2dW21JujhnhBCiDGqvVZu/CT7gZ5ximI0IsBg
TQ6h738zK/uY5th185rgE8alURanvC6BStba7DqgYIZ/v9UjKu4d1BTZ5bNuX/PlkJnlDTawgskk
xGbxGpWx9zuisBiak9Q9PNKkDoFKBQwAYKurdPu5Hlfs2ht0Ozv9AKrUFUHyiivIJJj0h6cbG7yR
jxRgXQosrzIAZ0VBVDHxDRSNd+vTMe85bKRlql2IeZhDzuuS9xg94nndi86aoih7MGmdy87axptE
kBqYHmfCFd4L5RUEJWm3MYsdCzdOAVsM6api8WAZEsGpjtjOpZPPoqmFLXdXCmOL++av3YIsak5A
YycF+jj381bf3oi5FHuJN46bcwHvzmgZRngwSCGzQmpF/Hq2sGLaQPtssnvEUSSkfeCAW6+FVYdi
eJin8/VEI5hJEuIr44A4VFg3xYx3HDCQDyMcf+q5K1O8+5IqFT0skQeddktWBxwd6rhrTdSEMoJh
sVl9KdL6yEq/xT7zOkaazC+MegLopmvhbQ3TL2FWLth2BC8YS76HvIqV9puRC+sqPoMsUYiloe6l
wnsJzhkEBzr5vUH63FZ3P7nMFuouJnG6vntopAw9QGiEx4phtVB7tZetg7AkEqBzdFOEglQasmi/
oL6wFX4wbBHcGm1v9daYrxnas2UPi/VUG2iSpseWRrvApa3PF1DFue62MybWDMI/iCESr4oRwMnR
FGk3Mxj9fpREUPqjv5iAIRkfxcw2FyD9oNjbMSfzMefJ+anNABaadMBWl0DJmH3N++43wFYGaPRJ
NTIbXIdZkA/KaQRoR3o/TegEC2/b8C5F6T+75Yt1vsvGvUoXhATU3WsLp3HSo3EVAAX8FoLuSDBx
6rOLOj6ZQpg4F0SCanHHsnqPYMVVfdLGk9Y+6wRQlZRQaAd2cN6jId8Yu1cLolmKXqdhjMlhS3Ne
fAMXp3rTg90Ddlxcf2TLnKX7GUPF+muXT+fW9PEpZMZZN0KuCPRsAuF1lWBFCfH2gikXPlFHi2m1
TGNGXZTMmaQlOfdhonZJsmjKfIefJhOy8pxbVCO5E/y1L8OxqjkKC0PTyua+lWRBbDUKCUTFJKsS
ArLi9VQjzzVfY7qT/nlU1i9E7gdWO73ST1gaOo+hLVSsCE+uGzc4uV4spEEFBQB9fgpmoaQa48wc
1LR9ICu477OFEu9JvTxSr5fi4PMg9ZOPOeotmKqxs7Lfru6oVWVlbVBXFmaknUx7jT0+13oGKyYm
Dqomyq0mhMR/vGANv674CMoX+UQMu1ow+6idM3vJdfjaB44B4M61AYBIJy05az+Q0FPt2sErVCor
okOgGOi8suVELpGtckTJVxvhch4j7d4TDgkDHCCDYLZgiPXmQgWqq85XN68wmohtVdcwyEnSHAwj
3tUldMgVmB/kwfRyr+kSwrR/74f78KjThApUW3+BOLbOW5OjY4G18oCi0b3Qv3PNiTfEn3zSeDc4
vEhj+xxNwSToRQlkovoU8ZtGZD1Lrl/+y3FB8R1KUZyHhq7OoLr1tCUgXTGOFXNP4M3Ulbov3VRC
YIw2dSxxs2adiR5l1NQfgmLAK+WoJ991xxETODDJiqTOAjQOyCEo8ingSyRrY5jVLZ/QvhUDJ5Kj
WodO+ipvqIoi+KaTmHDGxsgmB2ZQ61jID1kKOpyXSsgZJoxz9+6MNvEEyIBeCpw0wYIXGmz6aKsd
ERBgmqSRPe1+0U5OcOgpWi8nvJFD8rEIjcAA4xHTO9ThHxYfnWNopUoPx5pTc160etOfebziwuqP
ssTNVXo28XcOGrZrR9+UejNLH3ZQmZnvKxLEuvgeyVvSiFOMTtzUg7jeaNoBooZgAA4WZdtq3Q8M
ghekPv+gite4KCWATz2kXvyRLRQxm4ymj+O0NGF39jOf8MxRm2WKngbs35zNBQMbNzzzxyXhe4mk
eBmaAkav5adJmtOj818Or/hEn3KuK/qEa9O42a3gXw9vNDHhdL5a5Wl8rEb7w/SCMq279Pne0ZF1
qw3iiWONQ/zqf38B8JKoSGsEJaO6N4VMn4YcWvGzPKv7itGUl6aut7gZ9so9JrgiZVs8WTWI8K7K
j5hsIcLb56QcfdBpp1Ts6dGIothE2jfG6jQXTH86sZ7nd/I2Rt/0L/zW/cgYAE3bWZUKg2WTmZZ2
0AFvrejMLILfT+T6OnhvPv/4lZXy/Eqfpvm/7iNYMg1HBEuqcbFXuJ1gTRwb66zSAtkABJBb6OuA
H1VhQCOV5urGR4B53l3fbPwBddVf9w5rlVCwYXLmnMH9g1NO6x+V3sLC5RrjoMjQIIwq41Vd+WdM
/FGcyqLdSZEL6jU3YREtlglEc1iUMz7HwfSVnl+h+5rUC+wdRjKCx4JJKTnOaq957lYeD9mua9dS
07oRsriHmSMoBpjy0E1vswdqjb4Rm7UuGVv3AvuIrxdPvsZ3WvHvKXzAJC+D99VLtBfAl/Nx+2On
j364GLzGKmqLFj09szS5tq6EmV37k5L3JS79Qd+O51WdHAc1X0LutsK6ABXCyrGnh0gf2w6uHIUv
xz26uEi1z87WeeT/5+U/sGVoFWUsMBKDYqTAPIRZPjFVmhrDwA2nmByOx+Rq5fOJ0O9KMaIeuW5o
JXx8Q8VhYArm9JVD4uZjs0chVZQ6MsH6aEQStjuOEbm8f3ycaIBtdO+TsqfngTZCwaspxLcwmMBw
U7p3BTmQlnf/6bYrZLiZlz+u8bhXH0hz1ESPFBaz1hkStLQ7uiu7AL2FNoJj4W2TfRsv8rNV7Xjy
WjfwpiEPpEoyPFlBWllIo5rlZkO+fW9HYrxEHngK/ohL7/T6I9Hy+TpKfkqJNqsatzTmbX4/hhiY
80mEw1F1RsNvmzZEvECvOtXHU/3cJK+/obHPG9qtPWLu+idCwK2TvNlYgonMqAEqeCyjtv/HQ8+U
VVKFFNuCxm015x4s+pZdScKNaIWQN8QNTsSAfOoa5tdSgicX8pTr1jFd5cFX7eBASeS7dgLNGiQ6
xAlR91gneG7zSE/u9BqkW5/gTQDFy0s3hEV7LJccSXJaiPJnI32ROA7/WS0HkZtApvTrrqS8jVTV
pNfnA0yBDaSTmW69BzuZTZWHvFjklzlqDTCe0EAdU7XSh40hpIm4O2obNxlk5Y0sCbsVKrD5D7tH
Vt16Z7uGLNWFAelt2igiN55Kio2i1a1Y6pkYEiOhnqU0efBA0N+NIN2ZHt+xzbYgr0di45Fy5fKw
eG/5bYAQSPTomp9VBud58+Z5iZ2qGvwZ7HPUvctV6MoDg6sYgigWyms49OaI/AueOh48uxfvmA4U
jDZjhyksZ9PgmE/zVt49wUc6PUC+BMLTwjkQkyRFdtSxnDpTrdpvIiqkL/ZLOULBHL9KOZtZQecn
ZWmF9lQAGvu4qtsj3uJEjbiYzd+KBSo6jvq8k3uBAlNGvLCMrM067hcqtxstv7jbJ71fLLaSz3xy
nsnqDGLNYI9KeS0NnxRKm2F8XU1GobMDUoMq5W5u9c7JYSR12IZfmMv5bTLeUrggdBMn7qfAr73v
EPAU9eq4IyLYSLJHgvrceH0WREMWjgdHfD1gpGwigKIGVfSB0Im5XiDdOa0CX3zNMLgiXhTLIYpo
IBaJRPBGg3pPCIH0rYmZCSn9QhFnRY7KWCSNgWUKxesF2eSZVFTFbks4nEReCJ06S/6sSj4qUBim
kAk0pRgVpLU05BoYXooCO9QXX8Nkk9fEc44T/ckUUg4nRVx7Lu+qCmfqlcK/B45By4fZMZA6ptaY
gkcLJ8cH8mvE9yoGZ9dI6Rd/IrWo0WLF7oEpqr//vw6fIB2XCEGAvdXFn3ple0YcesYlguydomSc
Mb7RnKXXiX9Vdi9M/uUU+2/fjFGQgxedJv+Ckhh+o2EzYCWTCOd3KlHRfp60t2IChCpsGZan9upU
6/v3VVz8AUs7HgIi2nW6qYRCQ22TBcYIylGZUw5rr+jaHUQ5lVekTkupI7vbDZJ9ZERv5augLt4Z
ucZ+oWvdvWYEOBnw4kDGMeOAyBktSB2QNX7VNDXWj+U1dA9lLxaFOXjZH2zdwI3ZA+nJNHvjC5gE
MVO8R5JwVO0KAewZl23cLrNL8Ue5sLjkly4G7JH5lGaMTPxjIdNxl0pyp+teLCMIk3naLcHc5LVp
SOA3mplhqrHxHvAhZvtpyfZizO/ldIqV/7VW1sRoCnpZENpRIGYcYRo9acVCwIdNFUWfjluDWdyI
pSEIrJJx4iFsFcALGOOebRqn4zJLpvZas4fjTfehAuK8EdtxP8EJVlwAY5MkpJEFdeTCHCqQonCQ
d7W0dgr8nBB01uZKppc9sdSIuVOGWB8RSZN/5CPbjDmV9cwpDvugAY5+yyB+UItiWc6j9J7o8E80
CRXhPHdIwcmoOF0ppTxMl0V5eAziWDGTXixoD/UBOpaoo99b686jbrZ86GgGAvtYczX5kOuvGNJ2
sUWIx8D+HcOnuVBD3un0/RqwkgFBMvgn+CBz40JGsr691CtHF2z0G++cksjn9sRFoeBELrih02uF
tTZYxa54IrQ/UGXplkjtFdfertgR24UP1aoztKS1no/fCsWMhE+HletBTlILiEbGLbUzSwpFGPIb
fs64FNGsijJVHGsCm8tF5xPDtcHOjCsH9f1mdB6nbbA+w01Riwu/fH6djnaTeY6P1cR49hNuzTgK
iOcyLCfVCaVzynq6GVF/jZiqGylDuNYBzH7fCLqgwQmd5tLumrmHWjHCxJDzIXxDUVZZFDJPMBKC
Qmk7wNakVah+S41RrG54IEK6SFHi0M+VXGnxG1hraW7X5ihl6bVkrwEoWDgIowkDCN1r2CH/KOUS
4EBPUllcIoNJvckzdQMWD60lob9GoYjh/7iXMF+zhX8UnWBeZrQNQzlUBPrDyRuhp5r3gqGMfg8d
bS0EQOZh6Nk1RDeoVMw03cOGUu9+92D9wya4CtYEh/Vldnl9B4z/kBBpAv5zPLnobMBlfnx/14V4
aY8Rgy0vsGLJMpGcq6lKAT0FDFsPIHsYcl0eMn9a8SThEJ2ekdSY+NhtxxfCkS0chzN+T18mZaSI
12KiDjYi3tJFl1izJtvg5ctPGkjbspu6wWCDW627FtvWsLhjf00jKwDVUbS4qd485h+20NLZHYpo
/2spHzOlBVnAUPtvGnkLFtZXOQN7YEcQCdXocjuG7n+w/n/69JdnWX0eq0crvl4CSTW9ZGWk6aKb
1ZIDPNr77hr81nyOLt1hcPXa0A4qJqloK48aA++yccyF6mfugCdTP13fC0VbbC/39dW9WcNKWo5c
lJRTgU76F1vGPnd2+w8RV6KOiqEweoSd/8w39gwjVxVUkBBPtaUqIyzbVv7e/YeuNg1Zuhuv0YCX
OhugX1FlVwDdvUSff6DpjEUepD3Dv6YaI8JBlDoHAM5o4HdBuIALJPvG4d0teP92jdBXA46UuzAX
RJ3tFYUd4M016ITeXcGm2CLiQbW6xQtwixw33NjierT49kSBF89K3H+/697Z5C/nqxm8ciywfaaG
bWg8v1Dbq5Q+FOrgRZ5Vzjh8qYv/JPeyU+Tkc64eNA5sJtOyEAMXDlXkM3UqgEnElIRui4NEGbmn
WszXVpfaj+ECtExnu28Fjw6ccEnLzGEinrfLWrMO3+RD9MOUN3BsuhEq5AuJ6lEgcOTiDWhOz0AN
m2+bgEjOp6upPfk13Dk7TEk/jOEcyObpkl3ax2abuQhnqXuI/bMdXYGqEniXiUsyuQKVl8mTiq7s
hcNrVcTqr7eCNhiVMRVOcSoX16gYJ5z6g5GiRb6gvZJnn+baYPEfMIOBfc/xTcEnUNCu3nFFLeb+
0cSBOsc16xQkI0QIxxnSfqoQoZfCp0p5OGZJs/ONVt1p0nvL5EN8kuB/lteyq31XyTM4gVoaXRI7
uVjPsDaHjNfbiIBRxCUU9yWElse6YujvWsojR+xgxz2GW27vt8ICtxCyhkusH4tDRO2qoPKWGs+x
e3KEGnSFc1w4YzVdy0nFWOq1Yt0Vk+JV1EfrxlrkAlBthKSfjN4nr3R9tJw4Rnj7ZaizWxeBlp5q
CTmEzKeHrhlogLM8LfWmVHIVGWGQbmyuTyGJrD67UsIzFUyKxRnAW3RactGN/UoE2WLaK4FPxK/l
jziVoQh+fYfaIRKAnmuZgYRWilj7VeoTdCyL7cv6wSnYzJDH7cQcnS43JnXMRM2oV7lOJ0dpwYYU
sGWGCaPd1zEslfZTpaGNRsIq/Md/OGiDcRML8PEnNEIauargL1uJGGILNBqGxgiEwT4Swg6N5SHI
5qxeElt6fVaKJX9pVQvTNMEY/LOA5VDzBYdiQIQrR6SCKIhUtNKJb9c3HP+nEePseXam4CIS1GqU
jSvcSjJjQxsti14qV6eCiqvRRWZY8FH67r7I1TAO656GOaANRivJOAtfhHX8jPlt30WxYYJCC9mq
fA4nUlVDvBK0Q8mWr22zV+3W9+RWyJZT4LKiwlnp5TqAAK3KUQvWontviKkL9bGz8vtLQWc8fowv
rdS3jDEP3J95cFoq6RZGG9C3dteEKYc+vUh+xytk435Ju7k3ltg4kYoR29TZtiDFpoNqQfyNmF2q
3yXvjbLjBMzXn3YMYTjb79nKx6NCEVeM7shBITNJ0NMlwrM6ha/u+HsdDnhRhRaSfZKdWgrXqyie
A9Tiw7UpVnvUF5p9JRrFDcpVucnRimQvUkk4mwHWsOKz8RuV52t29h3fy0neVZkvt3CwwvHApQX1
1qIU1QjTksJg1scuwsV8vFW0wzQjLh8NgOj6Cegl+kNNx55/D+yH4abJhc4RSRKTEva0+oieyn/x
EKS0fVlXXd8D7vNSvE3a/EoVbJf0EQAyVHRvxbyZoYhOd+jyrIEo3H69gmBKsmjbkUEQa2MNqcxm
CRWfwUGI4y8/E1RcZk+U1re64K3DEO+sGWH5YOkww1eQ+UY2AT4J4l6loG9As5Pt/kAsI0nmPD1g
oytQyVtXDiV6wkU1oK74Uvg13He5EWjMNeXw+pPCnUdNhQnWTj+s1qtLABWF6rEnvPJeoc4/l8KK
JDgKwQjtWwo+wqZtnqjNfVkc9DAxmprFuIjMEU6lq2knaIAD8LU27mn2O/2uKNmi4SucItlL2xv2
aTdgr9orb4QSnQaMiGJypXjWxKpv9kcmI5VdITXnPodZjVlvknU2+CTu4Ce2giAEzRqtYNbca2C2
praiq+Fmbg1a00f/xxYdTlZKwbXEqQKtL7bCSoStpkGLCRvvFyjVhRKvXCblToMmDqsjKvR//TYB
cXqgPs0hl9Irr1GLQllZMhS/QdubEXXOZzzpwamcYc2mDw1QHRdVZZVd0d/7sxcgAMTxhguf81c0
UQweUvlJ1AI2P+kUKhh2EdfzgvbNRecpkvWRYKbTLZ1zUYmbArZiaLCsZeWztVePE/DcKc0Bg3f6
GHQKmYIBZJWMmzGMUB1ta/gF4fxjHhv6s6nU995Vz0dpQF72Bs+2NODEmvoPUoOD8QsioSlfUJBR
+QD8EEqZVC1ypTQka84ovwOauE2cg2che3vZn5BNqEqge8HCbDKpRWrypspGIvw4syIqUuUWSOg9
3rLuGe9k1IIw0Jlqm9HsDRJ84wQqa0IOTNavI2EMmKOtwufyGml5HY1aGLULfNmdD7Fx+8SmJV2Q
c89tpFkLBe+7CdagBzL0lJz9PKK79JqbK7G1CccIhCLcB0EoCAgkyHj8yEKrSC/07yT6fYYylwTR
XdQkPGLd5DceDGEZ1EKYLe77D2UBC6jtfKKZH2U47YNJAf3jZ9djHFHeRQTfK9PH68/CuBL/ywsf
I2dl2amjLfbmukcfzY2HN1pks/Nlh3Xc17Ipi9z/CIhzQPw6zweXfqiMRi3L869qY9byqDf8JuHA
YyxB8t1OySjBz3STVJLfGwYQWsv1D7oYrs4cZHegTc/Y8lylFzyEbP7EFIMq8SuFVskYTSXmGNmm
y3rstV2Ap6gLvA5045FmDyNEdNQeG5sULYDiZfvWZG1c0TTswgxuDMuJNuJ6a/iWdAmWIgR8Ht8s
niJPEQzHnem1rjR4HPNKAce1ixF9KIgMQcb6B154mlWZZAkj78+mT8GeRS1/0FQ07O/POLWoG88P
8b+/PbuX021gRgqyFovm+IMED3En1ymsSMfx+FVc2dnpBzY1UlYsuv9IOpcg4UgjleSLnGH4qQWO
XZr7U9EfR3kpImXS2YQ5C7Tzoa4ppIXBOSHVvpjIKD8ArQThiR1OGRowEp8Ch3NopsRX5cCTwLu7
ZRYvu37Js3rEHB0SoTv1NPwn74pK5ToQgQmvNaGgrN3l9UxgDIpfQMnnLrD7P62GufYlP8pAvpfp
ZEm2Y8lCGxIcK5K7nUy0oF5ShsF8OO8Lq+IDCVpMBnTO0yQpTmD+d7YQdLabWBOJ/W+eYQDKZW50
UE1URGFE2DeEYDmQ+NL5R0j1kye20Wpgl9HZslzOcHU+7bobt2CniK3YHSbqCCPC6wN2RQP4W379
9MC5LTPvq83Gbi7k6Lk29z/JLK2GeZAY32hY3ifmh7DpO5PPzOTWfKO+tXX4rbqqj4OqSHw3Hb6q
NDsdaMuePeX8bvSF8h1JdegvGyeUq5qwNbpLH7YlVB5XwVnLv+s5OJy6/r0vLAudK8Eh5rPe6FV/
ia1PTJ7mvJPxD2GkBDWpPKuCSPP7Nh7zI91p5I+meZgiJpX5VgRzMWwe5vGq1tXm9mcnmyY6dzZ6
HoT0FTRmvUgBgpTA+ai7s/v/qgXyvjb3Ae5A5d9IO7CWfoGM4XKnBxlpsrS8FgvCsRaxip1Yrlu4
7CHovXV5Ak2l/buPXAYtt5+AMD2cTUxUW2QnP9yYw1o++GdDF4U3miDlHK8xplKfSXnPTfTMTgdC
F7aDByDO1oOKr1f2fZ4uX/25qyLd4Pvdg5rOOWPPlRIEmadytArQm4d0Lo/lynsarxd7HbKENmuN
GH55ubkpjnJ/FseWGcDxWHRlIxvjnW/PJ3ns5Cv/xrdceoK66GmlgbGHMFf2VeAcunfOaixibiq4
dvlDF3dPwd5/GJbIVziHymxmpngeC1K/3sG6h1k4Au1YHl7E8w+p2U/QqhDamd1f9x+CRWsyzFSB
sjdlsQ83sM9K4t4g+CxXmAxk3UaEahbXqlLC16QjzxfJ4u+ePaMdO2SY5Wvq/oY+OlUtVe7sfAYP
ayuPq4UjBZXsGWPSWXPz2s98Lbj/6vCKCiclve66jlfN4IKLhuD0z8MblIWDl6DvvCYbB3wUssit
rpHuVDsrZ2mfMkadUD4ujrWdeN65hNs1Buo5T8sVqFxDvYtMexycJbeieEGu0QD9PI+z+rr/SvnM
fidVkHR7BR3IyEUHr7ekQiEjrBn8G8D1HI/H/O3em8M2mBwipMMQosrg9n52fBFb3I8AnriYhKm3
+O5VFxrVeOaH+tTFTbrFNCWktaOWDbumHI9mhEJjKvdWzdzlmCCDmMbCZVCJ0I4iokLqMux8tVNl
4FRxuigm3hKTUURD1Znc6mfZGkfkCkWldaCIsGgXZDbZDlrPcNV+uQJKSBFIJcwcPMOgcqzVukV4
CkdwpeRYKP1ETI11Czenk2+z9ELUG+LVrvhzlAFZl58stFuU7xHQamVt6afqbSKX9xw0T9+qvmcI
6XKpjhuplQjb784mKxW1eZHJtvIexWCN+HYW4f56EC4c4pWWENU9pOi8Cpm/X5OcE7zoCtmzSMKG
HNllKTfw2K/pAxhFjdBWskYk7twrTutjazJoYs9VdyItBuULRLVilxbwhlvVeilB+JGOObxXMEpx
lpMsQeVH8kDRBWaYStuAjKW6yO/Q3r0sp4ZFT6JB/ndk4IknsU688eJI8lxmtj4xBfoFoS6J7bsv
LVC4TZombMlXx7EhounCfhcomvusu7lMPJaTEA8sQo4Dd+yEKmoDBCZ+2gC12/78YO8KclpPjkbA
8CVeez6E2B+OVdLAP8VGcyxl6YBBjJIKCtzU6EM2/bXh+vtRcyW3hPuP4xcTS+IAcmsjxyVeYgA2
vU7gQgTvrcMlq9pjqijJKbMd3WCGUha39C0UkSwEfnD0YmuYnVa6G5+sq2s789hioMP5Er3Cguj1
CrYFdUBhXT7CygQnoBDCVu6xhAYdFaTQfNfg1D5qM4kyO8FtNLezhkmvR99R5b0dtFaOqN8MYyiN
3ZSoyrFimS0sLiLgtK8V5tielF6wUoOZrKJCGj7sXUYrAyw7Ew9ZnQUR01EBW0RgmCTUPu3nJdST
7iA3fQiXozIL/QA0YbV8GwnXhPBh38zcUAMAjh8jP/Zb31HMwi9tE5NBiCKbzWxxRn8D5602MdnT
4Xma6zIc3mUAcLBW1jxFEMogbZw82h5QFUsjKSrwKH8mF3gwb6CQmkLHRaW3EPfUSERTN8yliRwj
JIUCUDIpx3PwSiRpvlliUCraesKokas5tDumx8cB0DqEV4am1rPQCRYP0tMfe+1MnPD9S1giiPHm
wgJ4p2X1MLWYCbnNpptvhBmI8fAjlVxvMI9NHpwHSYbkItl3jYzmaexuuZntsXR5yCA1FBlMBeI7
zRko8jPrXNV6rCt6ENMGAQZrhxp0K0gXwTutm8NJmr9Dqmh/2+stchR8E9y+D8ny+x5MurHk+a34
swtjLzReQc3TMk4fklJ9jzhZLtyLLcr7/X2NBh19QTvAvFbImrq6fV7hHdsHh/DY67CXfEpFDYnf
spVs5i/t1mLMqxPzMs3c91pk7ppwVhtNsbX4I0/XkpaIVq8OOhUQ6daZWqqhUe7XLjyck1YXf7EL
NleqgjLrZl5sbeS13DsoAZ9yJHI/onj/gE64A1PagQJvH6FeKAkmv7l0OlXO4yD8elnHdrKVIKT+
OQLvH2Pghv7dERZLnaTDT5LIJyp9XPNIV/4TFlEGtAYqtOYpj6HiJm+ciV+P86lDnf6PjVUkdeyq
4hgfezE/oU4eMxhkHcfOvbBtJZXNODkJZMonRU9Q3JZ6HgTlAqya9ScCwblLoh/txG9EAQ2lImwl
93l9n8EEXi7Mc5Jkgah0prpPdImvb7LbD/oaaFV73A+NtyqJwUGlgRDOVFbj8/WxtBdjQVRY9xBb
BRqLQVBQO+GJTLrTvq6kUYuChk2dG4jMqQkzUKFjgg6xk5B6cexCR+pjsmAQViPj2wtpXX435xkS
0M5F9cHfWbSprt/mj6WJmUJiFnptjmXAjvPR53UKLxq9AT10o44OiYxzHNw6TY8eaECJ7u7LlMbH
QZxMu3bNpAJpqfpNcMo1mIw5NkWiFx/lrKScE9A2cgaNiQHgcbqtuqmuKmur7ZAzReN5x+Jfun91
+7L/S5XA78UH32VBCg3lGvSdU3cGDTvNKtl6QquNeYyHkTHZQFDwrqbqWnZ/vm27RUVR/aWDkkBU
Imnzt3REqh1U7rERoFZHQU5mQ2P1D6yV2A76YooAT6qa8T3bi4Rb8LM2ZBRCHEZ1F5u0jgLurIM0
kRqE8FKDN+BpTZuOYyEU3/+uAwbj5VwLIBBoO1nnMCxqYLHrBrh4gA4pFl/eZXkOfX+DlTTNq7H7
2euyGrBAhm5qPLAphTR420FZMZPFJi2JWTJqOzNZ4swfLB2rn0P2j8xVUKD+BWAWOFs9+ZVlYWF7
iJH0kE39ZqVaEzjgwVMtrUPuvYaDaLNEAbmrQmqMHSUeY3QhskNlFzNF+faHhBc2GVakCbLtW6Ls
iET6uJe4jXBFEtJmZ8ywIP9zIMhHnyesTWk0iOxhK9stiyr0d6SfnDnzbjo3gmDXr+CHB2TgLRDo
1zFooR+TdvlHRoQVxtXvTUlH3wgHO4EcJU31koJ5fEfkDsM0uGNd1k6BWExz+sXz5y4bAt9A8SmF
UNwLzKdrBcaffm/gVUa4ihi2RSLm6dWDpcqVHNdEaybMkki2oPKivnRgjPslunGLoX4FWKsxiz1s
d1o9tTgKM9a1puGPAprseiF1vjFFngnf9T1Q0S0gMvVc9ntBifxaCoLui77dELSUR6ELe8qKU4kl
5wQmcz7uMqDInW5w57OCT63wNyvi/RX3gztTyAntp/Hxixumwln4IwYDMJO04rbWG77MuDiIDhVb
BwjXgNFNM76YSBQ2GKZqeaOrNQfNJTFrLBE8vvNQPAflACShHIE+scirITPDS8depJuf4cRnuQlT
IQme7+HumWcU26RumGu2AS49GkmKOgWGmHriLGZQ183MgIwxwoORhZYuX3fE/VAvVqckBjxugvOU
XHn3Asr4yeV95eRBXWr4mOoXNcbIfasAurzX3IDfIdBeWEA8I4jw2yQqtdBHbeeMPc/f/ZRAoDQA
sBGO7/OQ7OaOPXL6YvEc7LkOsNl6hx4fOSj8xgjLdKaKTyGaiaNEfGCMpfv8j/XARud3pQ1Cfeay
NJtSbnyll7fGtAej8HbW1Vb8tqykSiAJgJhLj2SR6Mn/w2CTlg7RUSCTzIuofoBZ4vY0LLBCyWen
wOIyLss6mD7JqAX15Avt521/6ZCvTDVWep2qnE2lLKuuyRocTxO1Vzp1aGG/0sE7X4xqJ6mUWBIx
l/TDBERcJAWYJ1GsZlI3FZFoj4bbe2bOSOwFK74L5cw98ekXGH0G6NjKtTDUbW5BCJolldlAU1Qj
BZAZ+Sv41MSBQGpJuCsXE08iheoh4D5msG2D+MEaAccdBFpMa8Ct673dqriu6E5l0RCK4mhEjZK1
2JXgD4qxsbjxkOqUiZCPuaXRMuKpKpjHC0LJR6OOS3OGIVfBbLYZffo6ezOftIgIuZxrRA3RvvB9
ZrGBaYDVmCrt+rnitLQiOS4bq4Cl4WVtcgXjPzAd1n+GGp8itXLJccT+dqVDoypUtsbDPel5Kuds
mB0kdB0avhlgny9d4tO0zuee8d7ZZSJZjv4iUQfFR7OTBgWBX62o4/4Q/rjJPBhiElecw2sI3Gzi
cLr6l3cgGaZ+YZlprM0AVhxcn7LOzVg5vew4GB1+aByyYb8Rfv+gAWOiSHgpIadFE94d/ImapZpp
efbmM6rNshCz2mSC3rd4kuSfa0zhnMMq/Jyehhag0lORg0px/fmM5LR931KScGWzmWho6UhBpjxk
XjrIvpHcMoQ3pqgoZ5DpG7Zger8NOWafRBavSQqAXEfcQGOHMCrifMysD8KHtPMDG6QOu5MZ8iRv
Ohsn1H8tx9eGP1tYy9Iai+Je7onFjSjGqn6lpeD1EOzIgx+AApu+dQuAyhd+C536d1dKII6B2obF
Gs7Fn3SKAjaqb9aFRLi6fY7ZaACZk+gVV2VZz2J0zUnmCn98puSGeEYML4ToSm8sOFd36qdZOIts
PL2pPVvSEEpk1dzfHOExI4PBMSu/NKE4ug2hdfO2j/5vJyuvLJbjfxcnZC/fDS7CLqL4w7WhU5SF
+vqvOagkOMkFdl3L0iPsShg2vDuLCPRQWT5UkGGPVaEnV5JOhLmwhGyMjRTmZ4WkAft2Kdxn8VL/
sbMpei7A1SvgOVRcmrIznT9X5vhgsW5uXIEaeuOyZpbnRDdaXSMTektr8vear5Sl24yjyX+WG6Ag
KQ2imf36Sb3OlL7P7w3PSwWWsmzw4hIl12uYeS936umaARo/XP5Cy2xbM9E30mxOGVGuH5YpAaod
eK6gxerFymkYi4q64pvAlxbgrCYBW6y5QQHFUJrBC1Nw64a59ogOMvbRMKSY+fMFlvudvWkKNHt7
/1XlRC4FOMmIgsuAKaI9uyo1kE10YvcSzcpxeIMEBzem5KITsFeq1CxWJ/lFB0jUTdwec2gf1fSx
iTDiR9/GvVjrlecr2K7yKwoyF2FEavuiD2iQSdRI738UGiN3reokBlRmb4sJ25DU7uJQ+6ETJzyU
YRJL+nafindxPzqcj68PP1r7V9r5NXVj0El2nSFyCATFkfuTAKNWP0Xq0fqoVhxNrYZ6+NEwvlJg
z9eiDQFlwE664tJ45zBv5YMdv6ZwUw+YWMiDmsogTyocHSBzJTsa32y7SVfxg8jsRM0t/qQp8kri
XPYYuXa1ebfx0pHSAB21daVTiJeZg8pY36WkJqSyw4dx23ze+XWnGs+98D6oWqVNol5BBhH4UsmG
sqXd9LkxykZFUcXRUR1rqk4dNXXpzV/MIuESNtzGxxETUrTkDkB3OQ6D5ghZEDp0JHyFX4r62bMl
Ryd8PwmuVpaKz43kqs7WVea0lPEvBET0CeuUxUQ8IeXq6TAL/0L5YhQhAqwXssleRsN6RrQrfi3E
C3qT8P4MGScP//qNt7vkmlB0p23GlNJMwfZK9KxwBgKP5HP54tCOFcDyHPQw3hJIMC3f2KjMLlpF
mNgniPnH14MNMBz76F3JjS7sqKfzQ+QgZ1b3eYw/L3wLi5pAd51wAXdfR4aG58QR8FCdm9k0wCZE
I14ecopzfy0LXpB00KL21CATaJ+EdMKytc8XhTSYdhAVE/fRSfv1KAf9HZJSveXN8rMCKD92am0c
Yxh73Zng8jvGJbEEk3fCijrHKEcRnSgiIYll1GP8paUZ0Vl3nhtFxSVqTE8ERi2Ne8hevbxb8oQp
2uxL8D3ykm6Sa3lDM95D09n2/QC9KuP9V65tSfM+WQhMqH3cai12D6iYxr3+K+n1VBSKcJyHBnIu
BcwbhAgeUmS0cYPdOS5OZNe2Z9ppjMIrxsXJswwAumMjBdj44+JuBhNlb4AXmX0LRkQyMb8Fv2aX
4+aFv3xuy3GKFTO5gVlhenIvUfUz5LiTnR7pipB3DPsqGSKphUEu8nxG3DCn/FwlEusQYgZfrl7O
rsKa//sstAdpj6GB+0sx+x7h+V4DacpI1TQp+R1EIptbEs5NnpuSUAX8+vPiut7La7rX9UOGMP6u
UA5BhGOQb57q9+aM6gSIWgbwlO4Baniezs2utG4utKT00oruwQBuLvKDfANsAIyfgESHh7QXPdKU
N07u9sgkdF7AIMgNS2c/uIb1bpe1x9705SuDMTbQ245SaaMfBuy1ci+K3xP2HEKBzTgaKzcYWdlN
tYk2l3arlr+9rmX0RymyhY0xFqjvdv51UvUEXczYEsxj9w6ynb0Bnt83vc87G4Widv6mFUQ2m7sX
m044bpZkKtiVoB7eyb0Ogz+CQMO+qH8X0BrTXsDYiW2xWuqpMZKpzbwgY0ci5HyN4J4BH9+p4Rk5
zXXb9XaLKA6qNc9KZcCLzn6IMRKIfZeuEBuWxQ0ou8clqUqy/J+pQygoAOis3Zd+jyUVrsdI19IM
XSDBpOcGMVRar35KMRkr+q2/KOGP4N2jftbwFKWi3msjCxwAaylRKGOi0diTh0wMcGqvIQccoaWU
oGzaiMe51QEWJTpLl4SEKZwS9ggqZu+wGzawQXrvUKIAVZ9K50FkY14vQTn8MfbLEtuPkRgs3hrn
0jtPzFo6sQKFHaJ4JCmDMyNvMqGsqd9Xq9rmk995NKFvzQCB0PH8tlkdCSeGoqh5SDzf5F3C4Jc6
MGPZWZvld44U6/Fj3D6z1vYunTRzn1Wh7QJ9yIaS2cYDLu9x8IeQxgzYfZEjvW4Zn2FrBfHo+u7X
T7GZumNT00kn0cZZ8B8lwxrpPVjDbBHBu25ysIlTW4z18SMUd06TwkzHAv81yH4ZLsyhQb7IO/61
VnLbjmCoqHw7B4N3RgVj9qFSoGq18C+9ZDQQtCJz3YCFXgUXjt9HX5Pa+8L49UFvO5bAeT/PDo7/
xUUjvjaU2FqsvKQGMeZVnE0HA0Mq1/rsYFz18fgvHDlnHrdfMRtcGtfH6VFR73V/mCg7u2l6DrXu
umphgnDn3MMnp30d3OfPmdkG9Wm63xbbF2XjfPPsXNo/SuUo+n5MarDhBVMBSp3dmNKL43JwT2yy
uavvYDx8JsGBs8SZUtQRWPn5HvBRpxMENUOo9SGKsQt++RdQKw2Hwcxm/8iL4aGriYIiS0dIdQ8m
UuO8SCRbQn1CSfpss3Yhl953y4kFoxVVkeM3cz6PpwcZ0ygAG6ZOIhD1dj3BqxKm9wIqO69xR0xk
AdIhitcRE1NCaarZ0iGRuuCZpKsy7i1Jy/N0OONqQYnz6KLw7l6+KETytXtEQvQWVPDZt+8XWd6p
CTtafBJqJfCcJBs39It/WsRkRqg515d2G8rHQ18AjE5gY577Z4slqYZ5BIb/l4usYfo1M0nRGwcm
wvFj7BG06VMgtD27/YPMx5l0aU8kLxVRDN4T6QxvwmHuECi1GqR7B4ZhHaXj2LWp3pm4gshSEg8V
tOiWJIH4XTskZVckYpu/aJqptI+jz+8Nnqj3Cu18F9S0YVG6zJbPjkOCsV1EYTqTS2nCtLhCA7uw
SALWXTpnRC5GpZ9wbk98avYhkSJJL4cm8EagQZEtFM2JRFkjX4iXEruxNkJP68PPuceRISjjitZM
n7Yzp1HpdxvKx2jaZEyNZwESdtK56j7UvXmuS26M8BKhCipEM6V8HRs1uEPtMLgMo6rnBsNeLM/r
zRGd+hOtY4UpTE0IQZNIhgtOkmrnCGVSlYpv92TAUJAYcandY7nmxtBU0bmCEs7KlYTylJh4vgFy
3n4AOJcsXSHadgEmr4snCgB2ZuR1LO7ggChtmsPxpIh6/pgIOhEV1e3NwndRLmZ0SycIoA082TEJ
H6W6rVhHqJoqxcZzrF2K++VAyTP/dzGBLYy4M7gXq/vCFTCOU9PIEq3AOra8rQUI548AyVEvOops
GYbGdzrfa7hlglf33PdMLErd/tGuH47jDYVpzseGH9W5ntE+vdu+hPPlPAOGTBQracj4w6eyg3J4
w7TjYlVSrb/AWXIsPOzRIRKesLQUwYSRv7iRLzDLBjSzchQkXwQUCggsYi/o8IuJ/ViB8EvXD77F
151MAPQb2GRPAyDGEjKspABjAPKSY8U0Xm493yqw0Bw+HsXY/dAnn5wiBcQZGKgXmreRJahivy0H
NIveR/UjFvCDEokz06zqFlvPwOUDM1fIU/U6Dz7+xu0m5dPYVzKeu+3Xhkc+pE+pZAEtUELCHxeA
W96CoodW+fEhufs598yVjFGBHa2qpvJgpg5T8rUpzLXiBVMK7PSKTuOF5mZu/GKMUYLln0NLcKxd
oSiaWaL8HriYJTGhBR7QeHbQnx+Q3Y8FI4n4NCtImoB5dIlVBJRNIvfqtS9DSW8UvKlG73F9V0ap
k5V9YVyY9JHe30Bq8oHRXyZUfChJrazp85gegWr4drpOBT+yx+QX5B8zhhocRD0thc8J2YQSIpgq
0Fx9F95+wHEwqbUaQicFhFAUdnNI9xcorPv1+a+Og+geZJpyI+sX9reK5z6An8LS81DYlqA4clym
pU00ijq1aOvGn1AbwDAPmq+Q53RolfYGfmwglmsaSCs9BpKxiPn7Gyfn0NTlrix89OGDUf8fQCRN
hotlbgz/X8KtOuv20BlBkLxsUeQ8VfYYKgNWcCO7EUtKiVplIJsTdWjOlvtnQnRCUiqNz+uzcWw7
uwm1htzMKklVzUqOLUCTeWUoe0bVR18i1+gwmVa3Alyy5blExJ98ToK1gM9dTfvCMgbveIC3tMn+
w/i123DvrrMO7Jn8RteF6nFkuwnaPHBW9EuCOxueJBwL2AqwKVU8ZEp0P65mHP3DBe5tF6TVWoEo
dxNCW+BOYVXWRbfwK3DhNuaILfvUprUqcoHa06pRBIs/UNU+C3G2dA5cqbK89se3WS0NXRnDOust
kUxNF/enVugV5zPpWKMZfF1YYaoe8wgFqivHCnh6/PLhs3/UH44pCl3bf/zLPYXiWTamy5r5uAj4
6LY9GYsg/5TYBQC9WSjB4H/lCl0lkse9SaMrrNrCwm0njaIw4Kd0OML7kEe+h4CUmU9EZGhmCCfU
NvHwSKtQOzkZ56Iq9niYWgCEftqsuv8GAuGjSBX1ggQKK8T3tCQXUhbxkxw31Ig1jCwkb38cllZB
rgm8TPCAg9xBzV+IBCSpSp+Q7ZSqrQuK5MCj5OqV8xd+IemFWWPj1h/wmzJK+GqNMieaA+G/bSlD
wq6C8z1RExbIAkVXINV6ILFy5XIHSTBsfN4snqzW3p9FQzFAJ2wLf2oeP+eBIRQkP7owAqqM1VjM
KH5Z21cccznZPvfEa3BrhXoYEFRuSoF943kgmN73o8KSyBvSMl6jHbXgqonothgeAiQXQIb0Ltga
EsDNpuCTLOivex7517Wkb64RSSn2BjxMXJsVe2l+mtZDaz9uJWRTg1BH6nwbYYOl7Gx+/KYh8Olt
+MtPl6kWhMrNqnyQLJeNbnpyG+Z0X1AzkWcaxOK27eQ/FPJbhxZtj6xq/ug1w+XgyWvS990n+6H5
yO8ZR+o6Qc5bOCw8k95bujjyk/DSjw63Q5G7cotfTBCdZmED0L+7MwO7fc2ZnoooxUNCQ51VYFHz
S8qA2LNRQOZugnvUNcSKfMRucaWNrDDIA950e/VbKk4EJwtXUZpjEjOym1oW7woUWjPk93INBLlq
jfghSamU/fuf23A8lV7mZsAtAdSQGRIbMvnMmqh9Q/bFW8Nh6fmSDBoiW0Pk3UG5AKA2O9UC/Eu8
7ALST2vllDcSOWLmlodTn88Yn4tQXYzBFPi2hwUIsdLm8RPcQeXwlWLl2PXDpbW9HCTBQQdGz/86
IDbdiEVFFS77wQHhvZxsOQ1TEDnjF/zgMB2np8J0iwosFsDuWO3TfX19fAy3ygdfnviEtLX2NxOH
pIMWV0bwfRt0LC4V+NhaMARFFPS5ZwE+6C3517lJ+miG777JtTf2eO/A96ngL3bXZR+di9Xhnaf8
rJmXAWCaJbh55mlyjzk2jR2secLVPW2FHoM9zwT3uTjbglv+DxKyJ6vZgLXbz5KWcu8agCpW3hUI
c05tDKOgSAMEivBvpo+kOw5WwGvXmKf2cwKEhSeeQrXYVO9m+7U+eCiKj8SVuoABT/ECZNs3yy1H
OhSpK3eywKkm1/KpxOjn3gai/X+M+YSRardltYe8At93JdYMg1Bqh/ezVTLz2nX8z/Sm4C1ODcWh
4qHSz5GwFYDosGIoDwoV3DnkNJQU5JpJYrLC42OtdS6Kv1mv1aT04yzEIsTEsawf4U27bICHD+j5
wJsQWl5as7Ytr0mkcfnpSYpm2G6AgjgDSu9BlHeR9YsjunLzqF2xb4xAbOQoeyQgOp4BJV77Su5a
9DOkWOdR+C0aSUSP/5tQcP27TerHV/JW+ZE0JT5Z/FIQ+90OD1kZz+tNM3poC7DNsJPGm7NGDJpR
YBbrzDFmg3i1g14mmOzIAX+KX6kmHGlBBhAfnEQ9aEYs02JzKT6T5qbVedKiVBW38UMs8sILwE6I
CnJyHfQ8wctw0PDATjuAsvX0Bd9jvxchiZev8hmhO29sttAWbONh+LBcpW9zMLl5T4ZMjL/P8niK
OxvnWkIg4rdoMZw7LMKpl1e28QJr2mDrRMPKdRgwZ7yCacUDWx/wORPSdTxuIUTOgXo+LJH9O1hY
2PlWwdAXXaApvu0sJMq2qmTudJrBqew7hTHjnfS0RpUoPhpcHS3JOZ6fZsEFKZKmk4FhfJ4S4uPA
bvirLP/iNTVRIF66vDE7oE2c6e9bJ20De8+TipLGJ1NNjdqQvJmcsZLe0EB4roUJJIVpyzn5cERc
VvM2xGKb5w/+cwi5dK2U959B4zBTdvOnZGgjnyiCbUBqmQ/kzW8tsBaW1tM4HoOsNhNvtzpYIgkj
LodMH3B9Smo0sLwyTxFyYTOJCzFQPbqsodSTDI9StrgEcREZRwDa6dE2GIf6xMkVUUIpTjxu13W0
yL822meUNE0AGkJFA01mSpJMYDEYmon4gnWMMbiU285ZLKLbYkrRUKMLeFgAOEFBfQ8xm59Jvgie
jsiyRyvQovU7Fls36DCRpkCyJ0GD79hdO2Asf/I6LYC9QyzHl5VJQTLe/1rMF4C1SLT7T3NMZrcd
/5tibqQsAIXEAAKCa9s8EVB/ZpbsC7KI2C/Aw8diXQybscKjz1cJrhUsoqXoUi71PK1IVAGi4ZgO
ybYOnw3uVagcV+E7thTFqemHozhDfrNtViO1MlX/V4nqB6WKmBNZaf7YjQkBYT/8jrY/DzV92MY0
Wkl9m6DmIywsY6RoF28WXXVym2xN3uHqS/up6todz3LLXCTW7dK4CfwwgB6eBoYnYxvAFFeNJV6N
DpB+AczL+/FBZeqwph/+S9Fx44udT0SM6Dyzk/HPKhlY9+02IveRz1QkSlJIAzRhKkAWLEJvgr0O
2u+pIZH0Ib+V4C8b0NGJGq2Yf8pi+yOKWHSP86TNPw13k0/Lgc1AE382bx+lHVpEwiLwlsEVxrY2
MMYWb4Xja7o+36aAgL9kV8wZW9LL3bvDA5EEiLK2YtHhsx/y7PeLH3dMsep1MCDZn6QqPkPN+Ni3
AJnaECKKh1yTUqiPxKVDo4UKtG3PS5/HGB2sIuip1EuRzO1ok0xCicUePbtXP31LeSFr/n+f7YnQ
QHrCUbTcWL7IUq3LOLXvhv1D7Pe1mTv0odg83qp4gs5hPXInfulGA8Nz0RriqFRKlphNeJnXEwL1
HbZbeLHU2MMGaYSJsTPBgADi5rRcU/Byr3+ofVJl6qOCrkkfkzcovUXh3vcFBwUZgAmRcWgNGrkI
D4B2MvmZsDB1v4/PRXebx1bYScFl2OZFCa8wRdPnDmdlpYJBSEvQLrb+ZshHMTHoHg3PJ2njPDmf
ERvNsznpgb65VOJeNgx1Kq6iam1XP354ogTfhgHXBMwN/R3vAGVoA61TP+nF+j6dYEksgn2RlJTZ
KOCSaqKPaSXdMhVMJ4hVtDoyw6g+ldcko2qogXW4aTlZSPdnGfo6vNxPEaFJqXrRZTp///9ogxHW
bZ5E/TIEDOlhiggbtgoK/qcPUMVhBbZDx/n6eWdPu64m2BZVHWN9K8q/do62FCuUJUz2AGqYrBk4
fgPo+AHrTI+BMPTydxgQCVOYtxhljPn3xYpzmdZOnXxAmUAMsl0dqevF/j04XaAOIgjulSj2iL4h
WdQ77I6MdipVhx5tLbmN/3XIX0FggNd5B/dkfhYHfLGd7cfnjjxQjP9C3FUGdatbw+BEajOEHgFL
IdW1jZ2Pr5AYBd0FfoWJUPn/u6rjQsCjgM2oNeXs3889VmdAc9/hjRkgeZKJWg8hWjbAJrcCG6uj
0IkwLOJtXj7+S5daM1G1u/WBlgAbnomRsRr2pTUMqCHhcwFGrSN9RawV8z9LyolxIlPMoOjc6KxQ
K5FLYhOPWNebv1m3k1qM5x3nGOSq9frJRIqjKipM1ZVFz8IvW60o1SPZIE5Y27cowA04mgDGOFFS
1J14Q7jufRqETltdvzQsQDrYvRtTRtQWaCkN+tj+h+NGwB/KonLYNuPqLgSkv/Ia0SEO9GggFaW5
jNtzmu35i9JS5XlSNAuEb2nyG2McqpePEyAFVktHTLuqr/2+JV/hpPZMMmXhfT0L3OJF7HH8Q7We
G5Cx5jpjL3tB5nkTO+eXX8MeL3CTSZiJFZnLdhtS8T1Hi1Vu+lyWkU/xHUjDxbIn+um/LE5CS+s+
MWgs6XRm/55OLot2BmRW9KRT8Cg1jdgdZijuE0YW4RlGZ7zF30Juwl87/97ijwHUnys55OD8FHHh
XZsgO1QOXzHhnb+4/u+gzhxJGgfA4AOg+iClrStnrpMCsKcys8TJDUbYOvsJOl5J1TCf/2WPTMTQ
5oM2FTAfD0VqCTgpVCEwCZtD8b/KnvexcJY6kNuLhIRdKbO4CvQfgw7rm7gDqLT+iA7wv85OqxLE
pWEtIgtlfqmZTDfMQXtjdfBEp+S7UhIbcbiiq0pU1K83PCuJNWtVh/iuiN2X8DZwTVf1rgcVzZqt
hQTw9uaO+iGy9ablX0mZbY+XFHprSEb84wElmlEeXwV9I5tMDdqu76fbE/0Jwdi9Zlt+36/y+5NO
vNmH0lKx89SoUXbZnjU8NvB/KmN/hfJwOu1DasHJxBcAvt4tRQGlLT6/aHri1RhMZG866QAprvLN
ngp8pPfcgCIKgr0Z6n7+52CtRPMdmXmVD3+jmakZHPRyWjQR/ZlI5THoE2834Jtnl36Ze8U3GY82
cFgu/NvA3wDRda8puR3vF02xbyuutWnrcbvYdRRYmBqjFOPPYMuuc/WIANIcAwL3vMVkuDVI8fgd
LM+3n5Y//7pDWcqxFItczhKXTn3w7oi7vCKHTxRh6qoTqIjpQ3bhhXg1atVQtec/3+cUfQGc/7yx
ITdcBZ3tNFEE8ETEExdrLEPk6KMMmAelWOVGzzwmLtCgRx35/8/WB/DVLmOCoVXt3hU7SapmTLLU
8Q0ePIjyu+X5jOmV7Hrn2fvg9s469QxY1d9cAlCXzHJqL+ZzEiKRoYNX9qW+T8ajSq8nDrVH3W5I
YbvEAimKiTU4P47Y9V2RFkfNoLKakF28ITxMgTBcFuJ4Ec+gbn92Kh/LlpOlszjoTcKGppq04VZA
LdN2097Ecujn1dbYZf5wG5kHaZRamDwl4IYL9BfjZJNYi76GO2jMeHANzSSFgMcejKwHmC8MGFXH
BPIiEmngISERtexCRq2V9r12DQJwIFT7cTi8BDNPnzjNc943E0UjhWpUJLk4A9bHhh3mrntS02Y0
A4M2FnJMA00tHNQZyBahu4vM5R9CSmVhefPSwTF6dDx4gdqxYwqxofZzqfwMtKBt3pSw5dkV4Ot5
vUp/t11PFXqNHSwOYYf+DBboXk9hV494y6Cqtc+B2I+cgn6Q5phTPeTQ5YQpuPHbokBjaS8oRd7m
kSmPSsAMHYjIqWXPyUu30f9wamcS+SkHAb7bFrC5Bu3vS1mvwdLAgirL1g7y08LW5X3TmWkuJtfs
nc2cr1lrq8Hc4xRjBxk8i8tHGAdvr4Tr6faObXzu0nzeBOraqGMM9nC7AGmlR8vOx0VTbYu0oRal
65l6TyoHCANmYldDeiLFzxAzR6YIbhP3Q3DYsk+MPS56RDmhjfvL1WlbWq7zz/YXu2XdqBig2jr4
MuRuPJcE7DCi1iph+/NPqZ0zD4xnJEL5LEvAa2ntF+CGmbBxF9/nc0DOJZTNLkBYkij2b/pNFUPR
b3HWt1QhzLUSEIt0sSlERQ8NBPogagg71f/6GBfQiWp/H0wib3EqDkMe6eN8D5RHPuSnQxdZ2zjK
1fSw6Nqn0lW+7rVAAmNuwVo+c6Hlz60TPWPJSD8wr3Hxgum18fbcxmZ0Nv7/5mmDkVA+dGdvF/Na
4yxe964logxQ6W0qmF37MiK7zevPV+KedCeD9KxXhc+Mp4I9Jhh/aNFx5qx7ZdP6ik0F2yd8YehI
DCtIwynw3beJ3eEEvxN+o9XyJLDfOtjdiZp9LoH2/4AkRetxuUA5UOAe52GjV/o9tkCj47Jl4pAE
ZxSZcl2E+CONzj7zH/3jiNidP2loCBPeii0l8GJr3A4m3uuh2VCSvmFFYeZBiAAb/Gm7/tpZcBFH
XiqX3Lw1+h0E/YMnD7af7FpJqG+5OTSuSbtUnZiWqwsxaRDwkaz8HJtQA7erdlczuDKV3jFVICX+
KbUL4pQd466/pf1TLfSrRxYOyy3nM0uHD/iHelOGIXt6TVDBBZTYBtkQae5/4joRBaR+7rz/OiyL
yaHyiLO5kKmpqiNaGpvN48ualkfXmM4ZY0GOKzu8rIYQSbdRAevFqv3UZwA7uVXz5oIqGJDod12w
+THvFxIJFcDZf60R1BCLZaRDwuBVUxCCH8kzVkRE2Bgnadni5pAPHWhI+sZdnqHqzJiLv/b1zWh9
fmnIXSbYAjIKEjDG3BzCI5XT4P+7VWEC/UvUr5cdEwLeDbkg3K31AUloqUA5WGakAiJu4jKRkeQP
8D2G7ozjMdTfpy5FBOtZHh6vJAPk4tefnUIvL5LoH+m2Saw7uye/7/0N5/8unwUhR8YZNyeVHGgx
/vC6J+5kXgPMdL8HQ8KILXJTLSlE20E8hn6uYYfN5Y6sq+aSUaXFFqFxbUQsLdHgDI1aYsAQEI0K
aPHiZc/CmJfpTTsb/jxlCpkGPPfCyQUzTeWphd7nVwRSZFMQ88pYpUmw///S8YhHGQX3wa9niGbR
WbhIk5maTJtrO1snhkEHRG/yXftTb1orn8xtIxNusb0DhkBnmu8jVMXX1DBSEwqw+BS3chpzapas
CsCG6kWQGSyV5Cl2Q+egtpMFkYF8UZETmGUD+L8zrkfI57U5UJT70Y7lGzTruCqGywFjYuv4KBjw
8eljY5KfBc6ciGiAkvnimvj75xMhLuG5nXyaP9qUHYVP1wgPvOTlfvySDsdGFoedHCNGktpERW7Z
h0LFOw7JddXjzZ/95dK9BN6G0KrWjn2jLMWmCrZvBoOToIfBPxw7yDEcv7zhFXt0u1gNhBRd2F8Q
sn9MQx3lUADnUtOzK+wvOMK6ab44zRQRlBPnQ7k1c7y4XYoUAloPx/+5ITttbb/MKJt9XlwedXmF
jbLLTCWW/F/bwqaBQzxpjoDjlT+rysS9h4xqJdmX0b6MmVo1B+7MLLOAuSbRupXT2OMUnRYWzF3p
Pjdp0+yM3IBXX1R9vWlyesOyvNQGzyZBVgyTt5/aCyjJHVngEwQljDiE289Bq+WEJGEobSRCOgZ+
0n/XUNMEaWU5TqA2EcnvJWCGj26j33YwGsNACyzxm6zCvAuHXHAJwwm6n2uA2xy8CrGauybC2/Pv
KgANq0igTUxgl1gRe4wHL3LitS/rZjNouz7GZjZqTk0AJlR/+q7rB+FU0g6cNX9ghTJC5V7zTjkk
eHJ6Wsv6cBDugLsXgzHkG2hVnoVt3vWwqhrrbUEkyKh0XCkQfbfk2qDvnQi3W35PV9mlnrZ0PyE4
zDDoZtuBWFVUhnMW3m4ApeaHL7qGWqN/wdMcFAhn2J/haOfvZFCPGPbY/E0VqVR6SvNH1mAXxqLH
yX1hT8UyJiuEkOUQpSdU0ZRHSNZIdWYiWsBoJkW5dOHbZbPeRP83aRAPAAgQq2BhUYlKeiSmpWAG
pBFxAdR86B8+rvx2THFWxJaHBqWR+o7I83JvpbeKEBSPkNp1uuQipgX3d/o52p1MFTx980WrKnbI
1dV8C2r7EGUU+k/T9uVnIdY/C/MeTs99Kb5QVFQ1L+D2ZY8asXGOVsrn1Zpg0DOz1wPeFr2ZL47C
Vp0O5wIUrVXYefbWbjSNyyqRzh98SM31T6hv/9XW7PTw+K8w9Hwsg5vFUXxvkm03kwbDPrdv0O71
fubEc0z9umX+k6CtWB8vpxDczQ0tXK81S1YuR1M56wnYQ4zNxOisQyt4Knacu6JZbbe4CmCc4P9o
BA8Br52O3EeculdOrSWspXlU4XaaG1w20wLLIgmZ+Pfl39J85+gjRjCfA/U52NRwRI/Bq9LjtRge
kvVjr/UyHH7OsPoFfBFgW6PbmGr7cjUpJ2fjJrB7nC0LbpFlYkkSeHgqh55YHfqL05IE80bvpaLa
x9hoOXit2vdatMPUqNJgNT3Y5DTMNeL0+8JXh0W9XfHjnewuHyxwlfoxjcvOhmCjbNMwNrMQVMUu
t1S+t7Nx8vtQcI4Bu8jP0CLh5HdDjDfLEeqlzhQzZeKYb314oPwx9oEykgVhGfvyqCjZsduYqmO4
jMJM+BA0xg0XS/fTakcsM88Dq3CgH38pm54f4ROO1NPj8WTDJ8qFZXxzysr6IudNS+pSt88RSa+4
uBnVQAuobAaARIx8qT0i/OHBC/HPp0ZVpjSTNhg3VI43OoGmxeK+J5qRMFLCz4Un8hrDhNFGaXAs
mDj+lE8kBds1D2Hp7kujY3R9UE17PpH3gGPqz/iroZwPnRxsTSpHg9lizfeSxAkg8WlTikINQ6rd
oN+N+JY4UeVbMhyN2qnQOuKgcSQwZB5V2bjtjqlEFYEXjZ+BoeVgf41jHY9DixWVybtHkKk9As0o
Ks7SH1BfyKZEspO14AGHsNY9L7DW51e+mLExAyxsv5Q25hB+3XQEsi2WsNxrCvui1b88/2Mlpl4K
5tyr6/SvXzs0uMawkXEetM28YQDh/IzchEQcAwNr/wcT23BHcG8yL3tZVy/PvKhzrV0q28R3SqbB
r7eIvWAjf8D1GEE67QdJaago7UAA3/fwYBMIer5VG1yBBngOR7bE0e01mSj2y4eHG2SUg7oHo8sS
1Qvz+7UB0ERpkarRuNuzKeNB5OAh4/M3Gm24VdWyDh/dLMTq8oVXpvhUR9eSntB3ldBNJfokdXBF
9OdLlIJUFIJkC2CO+lDnTDwKch0jDJeeag/NZi1aVUTy9JZNaYyyItRVvnZiJsjMKW+cWt4i2ubg
F1fch8c+/R66r1+YnsDUyeEv/IEaMoTwuclWXvFbqr9qP1AbDLWPqcVIiLy3Q3grm4hL8yjk2jSz
zzsoEEKcZINgZrVsNVO/fr+0yD7jjU0ul2HK13g/syHXMnGfjMV15MbQH8jrJXpMC3XgH4mmnsl3
60nzqrG9Hj9wxCzGI5Jgkrxl/cb6Lu/FHhhpGlHlxQd0A+HFfMp3rRH0URsCuo2d9t6QAE1BIeOT
Xz1l4h/CReGJRUKE2bNTSjxS1urzyUEjhHq4aTalj2Xz60BBoWP0yKMjHfN1LJQbydTMugR1AE7i
sulgU869G4YQvBLJuA8U+37uN9Y4UwCATmCmtuve1zAFrwsdwgp4qzifyzsO+T6ZAkub/5salJHr
fQCrrR36DLVE2+mKQzxtv2A8VAvxY2tKg26/zfEF7Nt1wwEQwUPvB/KOci72fOeBsKTfZEXCSB42
Nc6vnG4psvahubKLubyIBFPwG7OaDbEaRRftoAM/0Gpb97ABEBCCLqOwMwhlaQnK2upTeud/9oFZ
vZpX7cxn5Azb2voN8u/C4BeQXJPmpqHYOQTaiGQTMNWzaQrXcA0GOgsBR4ZY0mNwZNa/TPA78309
WyGcJJPYRgmS+Q600PLGTqfvjMPUt1i1ZBx6f2sBQwXIvCcXZyfCJ5V9GZ9ES0zVOcH0UQPTlS4u
ojIBqVE2IQt7s1BaXvc1GabdMz2LaCkaleAgiQdMNlJ3U3hpWwtDVpoHHFGOipSc4ih2CQM4M/lm
pyuLrDRimIYR7gANej0zSOb5+59I6TxGw96cbzuKYXGbZIJrG+2nOAx4ZIXIPkqM1dfbWvaSD6FT
l+wY3LrSTNz6e0edFaUMdByokPHjwzN7uf9GvAIdlNIk9E3o4uIZd3pOcuKriIIHtLmbJgkfJYFP
3lOisM9ThBu2E9OssvKSLvZB44Olwihu66Ufy6DAU5nlJyxn4wxyk3TW6vig1Q6cyfBZQXk4FsPP
yH/JWZWKCeUOxQ+0SMROf+CgwVJlvARKx+FnwveRqq1aIeScACqqutQy2e+o3rLf3OqQCxmVnEl8
Xs5+btufbRgpnOmtmNG8D1p4I6PnDHCJXruhIuoYzfV3iQL4bxeMv/RFm5mqS/8GLM489hViNzHm
djJdBZ+IFQW5qeKcqr8pdsPqSznU5vFBpT/pbHdPZ4LRcnG9miMUGOSRJMZ4HFH9BCgTX8iQ/o0W
60IineYclz0yu2MfNxMsJgEsmtyhH6ALNzejQItrIF1CHXjNsF5kNtksW7ZavhWEjJ/msoHJuI+e
5sJjoUGZ4ukK7ckhjmZspKxQ7RwOPV7MQ/VB1RyFIxL0qX7AW0CaT5iW7bD3bFrCBnLWkok9XwQQ
t3pXCeU6BnmqDtzkUqOyxDgWIUMTtoVB2x6KsdlydoA1cGDwZArO1wWgBspDIfJN3YxwXci4cQ/2
sf9pxaKAg2bie81n3L1sfhbHKIjCkOgsi3wFjbkf0J4Oyx97zYM9eOUdvsZyRnixQf0tECtS0ZB3
fZKr5TRN+ACfZ6jPe2uu+dZ9seoGkNTpo8aWvi3e+Go06dr21FG1452BF3osXXTvKJPvqqEdR9LX
0O2g++jJ5gUWbbI1OVJThngCkzbrHNUipc+BFL2qJ2QXicmIYtHlwJ517K2/nI+ZKcUn2eww5C7z
bun5fHVo6kVC0We16RRErev060rSsNhTSXfZXWJ8+yC+WaMfguUj2/djMaB4nxuWKCwRlxuP80Rq
6ol3GosSOAPMWwtZ+EjLHnqNnVCt7LznVwGu3dWyE8rYjrRxnbjfJwEvKxd2oQPnf+3iUSlmx/Bk
vEwGb8xHi8W9Oipl8KoQkrBB5KpKouC3ihqMXljNgesFQw4WWMOS/SdKyZmWMnjVfI9DvWu4f/WV
Nm2YFb56BwcEj3CmWtjSGVME8Uxz7S8ksqNgK/tFZ3J5Bd2jWXDLy6DAdL8k2h1l5PWpx2Z6bkom
VixfRbAPjVrkSJ2N+bSVUT5ZU9AENTav+qh5VUPvNSx8XVtVqTQXVAcuUQEmnuEErjuL3/K7jgF7
hd77CZ2Qb6CBu6UzguHA+yjCQFmOk0jJ/ELKzgbMmKePcPbENf/7i/NWzMvukcbm5jjeK9H+qMQR
7Zkp/nozkNO30QVKBKU25+pYtGHPF1uagPYZkWh6oq9BVW7ovrJSzLF25TEVY922ZGYXEZ+mgUj9
Sco8yYD7+///rUTW2yZgjFkxDwXoREY4Ljqy7U+LNJaHtVSzoWxGrZu6MnCzM17MSTXsDnH7Py2X
ipa29F87/qgrFz6V3NkU0NmqW3uhdAEgfelC0QSyDaWcZEZfMaQtq7HiGndTOSRXasdufPTbhf6v
6gDmjL9EaH77wDze/UnFmLIFAjaXyhjz8fLTC1Rd23S5ihTgA5qwa3KHvCmI3te58a4N16RqNp01
Dh63SUsTP76N+IPxJWzZEhhC8vHCc3c+rCbTw1zK8Iuek2dTPEjig/qGue4JzPq0how+3QU0nMZb
GfXU4dY45dX8O2Fco2DiPQ5uUuzkTa345r+aKu31EV/qMb57zJkCHX0mOe1nm+q7BAMRQMx+hWPs
Ynefv8hO1g+DlPWtkl/xS8T4MkRMf8hVJ+raPHrtPlYGHscpxW4sOZ+No++trFTmYxKRnpucRL62
a6kCeKAFBilN+h1nWFctTH8BzLFAiO1uLV3oltVuBtkEiWKr8gDZsAkeedgaAAIIYGHv85c6rcyD
vXUCSfQXEFQcaIHfdxq+i+44eImnBmJfgpM9yoMdQFwPZS3Ps1wMHRuWuZhAtWci2kaB/Xvce2AP
KQC9pKMDDYGwtetwKkWmNkUNOmnNQ1OItrwGqTHpkBy1UVrLlIVjjxvovcwa2DxbgNeOHv0enE1i
iC/FGBaUUr2Z4OeGndAmxtnXsqi0he3IxLuosXKdeonkW+OhnRPHGf8v/N3FaL64yMyz/mp1ksOO
tZtvq+7RLJI+SQfADHT3niO69qt4tCPVwGDFCX2ZCjdrp2mjxqKwmK2106j5lvMgn33ual8NWq+R
1SIgrbHYz/qoa/QB6wvfqPNKYA0WVQoLkntLJ2XM1T6YHpN6YmmHYDVfzewYxYDwKxHe//xMClRW
8t5FuSeZa8e/L/nCkLtY27jl3C0M+VvJOIbbWq0t8z7HnQSXLB8Lvr4e/gDxs0ReHfzK+SDUv/im
BExzlBzyfU7wzlsS1PjptPTBnnQjUQxOhMc56PQHeirkl6xMImx8wgStRVl42HYQXrcbqxCiuZF4
u4vQ0eCkIvcoHOkNmqktW0G3gool97JnATvYQWAWUvctUV2dtDhBrZeD15ROYnSXYPifP3pC+SNK
IDYv+e/9JZ0sdPLNhloSucve5qkMP6vLcd6ggITfDflYA2S8Q8NWeUUMTBsIi/IGsO4ZSei/rx10
d79J535jsqaDVutmsiu9xmfVhi7xNOw26m4mfHEA2TSn+qFnuPLgEpHDTPgls5AkhPlfy+ixDH4I
zWT8n4Rn4A3zjSivhOJHqIOWk9YUImyGZQkZ240aEvV5F292byeFh/9aWXFjY3Al9FoWeropGYPL
NxodGXKfknYqPXzf0osGavTYCOIhTCX56yEcVRjyHqWrlvA7wT9SYhQ23bzcHe+8kqYJSGvjb8tr
dixfQVQeRPobLjYYdFEKJuOIETDXgtf0dsvMX5HafLgxt5p9Ow/wqgH+AZ2RSJUu/Z85Mvv0dONu
8H8iDLOodR1tjcXMER6BFmH2IQVhIu9yiSRw1D6yujmItzd1cC8dp0VTYuKz8xRULKZsul2eiX8t
KFvnNlJ/lPZT/A+RamPXclKH+HD2U0oiK8sYhDRVIt2v0TUxclR1HkdmmBtZcl9rhVMpV1eUizYn
S7fk45XR/n95+tDaX7aS+k/9wdef694Nf+i8EhBoRPT9zYVIX3tZgM6/IIyN0TVEOeoQytXbpHS8
rTfCeCrtv1qqClArR22EmCE8YeJiDH5TJ7NqP+2rxi7yw5ERIp6BJzCGi3GgLv+3A2g6vIPLcaiC
3ugJQOTcu5NdKaMTMnL4HKkP/HLSEExc4diU3SYz1cvZsPrfXy9XeQP4/ImqYTMhkGKNx3tvs6Hx
4rHXIGEhS8XIw+TL66Wjx9HJ0lPf3/wbw1FtWOUJ8ldkgmcJY4Yo//cfFlAWB1LO1qxahdUyIvzX
ciw9cJiWBIXDB0LdF4S0HDtFX6Do/PXAJ0c4fXZ7mowq1WklMcDPbJNrSR9fkZ8tHgZpziKzOJ2j
y1eOzunmTy+9ibJC5huDjEbvLCg39qAVjZkoByOsFpRbKt+EalYU/f0Wmq53mpNDKrV4T7CqZCU3
yy21eQaML3Qcw43I3k/lYWT+TOGxYlYDtGb4Q94wQCGay4GcSEoOp74NuMOLIlMNdQ2iYukJZpAr
VA3Qrf8umvm27Cg41Kd3LbUnAmdSRTErL0uoZ1jpuMrr1FTGmn/kXAb/RPY0HKyi1GJ5Yp3wTbWy
VluG/Gjtu+GTP4X8GYBVS7+CzKu0OAxsMw6W9Cw4keOjb+yOiZkmEzTjsVKRX+WOzMXQ589EgNC7
OSti9RB9WgU535uFOz5hmyur3+0qgs+Zqx1F4mO0Sdcbg6a0u8AOz3Fhcm15/dgUjbki483at98h
0qm0UhIzeXmUcxFKx7fOFVTjTSxnprFrrHVB4XRKtqVVuhQvOm5D0MTjvi6WtPRQGa1wZny/MR+b
0U9EDMWL+gp/4sxfCkYR2eI5U8/bGx8QzcR/jhUSs8Ln+G58/X1/B9wPiACLHMyQoawrOUJ5gmfC
yI9BA8o92Fws6Xuc3byVjZONTUD3hYwwn1ge2K5oes2NFR7K8B5wDsoDKFqEkSvCu+gqGS3l84mk
QeKMY2XWKSa3oSyd6tdLCwrwEdGu4HIThWtg0RpHYCjMmpLXp9hnAQQCfQ0EkTAyCR3dZF1qULNJ
37B6bib4j39Dk2cGqyBDFBR+nsdUyk3h7PY0kq1EH7m73IBxOJV9nrE5MGEzqWwBx3aCVRxBgDcx
6GhfXZ8NLyNl1jJ39KZh1J3a0N8GBEGKF5XE65JSYG3/T+DcW96dfgD1vwFNjN3ojoLjqQ3IpKDi
g0cl5BhuLPr6z2L6Q6fStdFEeVuWnbxpJMF9X64Iny5sYe5BK6O6Vs8FUx5b5g9JcYB9TGKf2HlN
mypC6aSIEcJXEvtAbilAicFJQ2SwIp0378NSKoMLdelqsOPxA81t4qyiQHdBk+MPtNBVQoWS0V0f
bkxDMXqo7LTjbEEDnEYUpSEQxA/flOrFPevqCRoEisUMCrZBokpH7S8tBuhtYTZAm1HVpME3OtCw
imASfxJuYjiRV1j/UdxgcHCtLMRo0IRx9wK1eTYaZum5JI5TJ+O6zJCHK5e5iRe7WowDRjH3cav0
BbmCUDlqIp2s8vueBTANdpn9Xc7aJr7cOso+pYIUG8DEmDJpJYp/WnlSObtdae3QanO4uDZI6D1R
sxeOZHx0UKowrXrD8/xA7AvfLXxlHMEUyEPE0OuVpWoqaJLORpi8O3hJRr8voKcvBDGF5RDEgnkM
yjFqKQjMSWPK7lRCUHKBo2H8s/fdzFvfi00ElaufV1TaXR897/PvTfkFM0aB0vwgiMEjqBbC1KSb
M/QOqWgBrNGdlEHwXSjEodp868fdN/Teft+ru6g7oRdJYEykPr6iO5lrmAgwMrxYuFH7qPL9Y/bI
pnswFDk1ciV11X3kbtubN48gSWVzQc84M7O+XBc1t8jUcR6kPiA33xGHjehInaZ3Y/lRPBgafQrV
p6uQTgHBC1dbmX1wr4zhSojnEVCyKDiMQ4jCYYNNybwX0uyaSd4dkNDKKQu7PiVmfTPNXh5Bnjky
mjnG8IfoD5fRHGIzzj1I3I8qHQOLiHA2QfkkOzDcQc+kPlmcrCIuhNRQy3q2leAQmOlT/YQVj7MU
2IZHrEIwVAEA46b7Cnme5gwWX54T1p0ejDvualKbE0pFhxCxIGOS7xoTF62lpBAwnTb1v2okUUqz
lfLs0rD0T0E4eGf4WMBA3sLybQ+wGPnGC8acVxyV2W6Ln3scPC9zkEjndbrFWb8Xa0KD7i1OHpNp
uCEkJzAHCSXvhR+Cixzq3ZKEhiZSuLyfk9gG/LZrqBqolodUqcqb1bfpsaFEOLjV6jzWjg8KAq32
X2TVC1ZsDH1N5kZxeXAm/cE4ZvhrVNjCynKQS01ci+pfAMPKqVzi4qk7Bj3VQjagEcQ6aotdW+NN
TfKIIYc4hSUTQPOw8InzTu2gggr1Ob24D6rPEscaKjxLchJijF4BBfnPXf4G0oLqTU5MtiwqyTBz
x0lO9w1nwdr0TQnTDuf5QhZCFAf1oi4EG1uSqiew6tCBj1RLymMqMJdQjfVZJUl4BnlyVH4m0xGT
eZsAMKDC48I/zudlow1dtIQAt5sY4Yf8lt8Q+BP0AHt49QgP6Qg29vkzDzyOgkTV6/IDMVj6NOML
YuQD+dTA8fX18lyvAqBoR6rEt8K243qioZDoADlcK7cPefl7X4rsdE/s5R9LjFYo0DEhrv0b2DVy
unueHwmfkSBfGMH/2RR7umINT0o5epUX02fwwLZZByNUUFj2O4wcpwAfM9jq7YwwX/AYLnguOkIg
NLu631vlHysUJ5qDid6BsJFH2uzdSZYPyOoHo350KC9MuoVAm7FrtCkq/vuqRRVXG+FwmagTQI9t
HB/eS9iQRjzWrSNGXFZ/ZI/INCbV09CoiVXUW0cSdDw0Fhuv8yUNaruEeOo8ui9MrmfOAZYhrX9a
C7wbRVl9N7bTjFw4F8dWI8/b8qjnXyTjEqttJajD02JwtP1RgPdenhdFL9mg/nT/FTSXrnmzScWJ
pCzrPWauROWX4lMvg4F7tfqXLNfFkO9UH+bTCsF9+mWJoTVU2oPuvrpZ2W0QrxOR0S3aW2dfUQbu
UfLze0Vdf4cHeQEJx6QbpfHLh6CLOrJxjtiPySd56LFBRWZ9FH8eh5IubbpNsd0P9tG/AEbZagYZ
QzNL70iNwMI7Ay6DDBjMYsfJsow0npX1Nu7adzsedyIpXi2ANR58qQs6VMGSVdI/PuBPTMp6RNLl
x3gurHZORFbFykVIEbjIPS9NltjKhGUXC5h2qtQcrZ6UTWoTBSsve+T3x24DajtVewoNVRhMHK/W
WoBCvMyTAfHykhyWCSBpokeSCxlvjSVwBtCcic3yzXVakTdDAkwsc5cTVH2GyYBRIkptSuHiusAh
CNJPDQwfoLqxi1ePxXtBm8SdwALafMh7eoWbEC+e+NWv+CBK+y4uk5Wa3Rj9AnyQS3SaZgUITOgb
59Uv2wmBkFvqmCm10NFY3XuAQopaV+2zry9boZ8Tac2ZRzrsx2huowOfIPxydbzuFKuq0Ff1/2bq
PWlC4Djzl1uLp4pWyZ1Hl1hcdBb5T27T1Veqn9I0hJ7ridqgGU6TzL1grGsywYunyru7yz/CwDI3
8Lt/rWCS94B9prYQQR5mR6aeC+WUzBetncmlTFZ/3lMCewnl6PcSVCzQd7lfp/CzdAV9smw1zbfH
YOuDFD0ZLU2xf3kLAGX4v4ytx97tORABih/9scxCUDgVQ6GhXpNjvA0/r5WSilCVH9tmKmDK7Akt
4B/QHQ5Fm60kSAYjwsrSGICrFk3D2mVrWFjurxbjiN74t8+4WSTq+oTM1IdSWith8iMWXJHqeLX7
cePHbTyUOq0Im71Qm7RvZZlXblqtgHJDe2hwQ4j7/1W2jIVJH4CgdBvvIfQ+N+LsVXdUhy5L8x0o
OccVhtJA5xq/rnbH39VXtNujdlh5hG/mTZditHyxRSCi1IWwO5rTT743j6SkLUIbPy6c7Nc2IdaE
nISaSHYdAEY4hga3AEQWP7Fg+TfRiiIhc/P3yBztNDsm8nU8xHBCbWQNK12CrwZHTX7/OhY0IJ9j
cp/Q7WL4ObLZ2/Eo3uE31aV04eF7YDOP0GLVUxadhVGp3Z8QC8sjlf/CwwkKM+xYRAEj8eCNtewf
WeWj4a4q4adpFEDK+NkoZEobgGDB9/0nHMxW4McaPVOGr6I3sLNOxqOG5d0ZxMdkDC9WyujNCV13
qGzB6h5hcKmNmZO8PrxDTDk047zRm1TkLJOXLJmDNaOuTqNwbZaH0RlHM6aNcrwuXwGOXUKy1gAY
X7S+ewb6cHcpv/vF6ZRs9qFw+xeP3IjwGcvBlAzHfJXgMn7aRdD8758pPjRqw1bLPmD9+z9dlKrd
P5cQF147/GqGFS5+rjO/JFoTgP+IOYrpgPOTgQoep9bQ4BPXRZQo9/9/qtmcSs1t4nUwY7LJWQQ6
xiC2USa3ir7UyzvyviQzfkh8NZwQPbn9dAr55OZObGwXw6MRMSgb7lxfaamTRBtHBKj/z5t0ZyM2
qb5xO+QBH41VtlSvy4yHRYglpHLFMUeitqGIekYLtK1vseF/cBBdmO3s/SbXWCczK9ubO+vTyxBV
qt6JleJ15vLYR5aR0dzPRMtq7xmB3Dj5pxnh9Ct7VZiC8gYTDx4dffELDo8dJWnOnvjgVPJ4DAca
9R6w601sApUbSxTIIu4uKuWRDMmPSP1DPCZUqFJtjEbn/EhzNuH2wc35fN0SFHtQdev5I6OpNNqL
qh480CR2dNo+VXbY5M9IprRLlsavnb1CMs+XVKWwuGZekDeSa4RRyDu4QQN03yDPyZUp5Sln/Eu0
hYw8qFTPazW5ODyZrxJB0mgKgS4OPkTY9I9oIpO4OClcm5mq3Z4uN67Vi0bjJwerxClCHwvLsJUl
YszxHJNgOPrYwgWtOQxmw1+r3fVHLfg3xKnBrwtz3nR2h9fB+D2ANVby8GIE0S2ZUezG1d1x8S4d
u5OEdoqMXlMAcRUcS8jOTCd/46vbBMsOWDLyR6b70OkOIBFnRGjN7iiPsNu5lc3KeejrAutOfAkq
4jxpMiPhHq3OWpUELOJomZSXQ170vpxyFpq6WVni7ALq/JtdILU8xn5dSDxDhTvX6Xk+hEAvXUPe
eiY2FIodE22ZdSu/FJrRxaFzMNvuUzyFSSAAnOMlWQQrAVM/vAxE2p2PQOlfcp5GRr4kcqjOccnz
/7rQ5HjvhwQzn2HbMZzzsU8NvW2ildf3mvkc2ChnWF+BeogSJ+lm4F2S7fIZB64/YXTdLQlT6LxO
qpnZM/WTL25IWQ+LX3XN+C8ROGcCY9bLJz4/9J5dX77WXCNKepkkKVDyGIJIT/a0kro5aonY5Fa6
UPqqzw6OZGTlgYc73tEtv2m+51OfM/UDazrUnjB2YKZ/Q6lMqAQ4kW9Ay9cgLyh3s/3MKWVaLvxW
hntRU9kbShktXjN8BiI2bSB376wqbp6vjfbmBMRqwXt5VX+n2f8gwQ9rd2Dpeny6zZ8Wk1Gb0ZJI
vNEwYDDrhfUnVJy0ElLlcv7y3XNvMwRgIUBupE42FH2fn+uaSNzGQotv7wzHkPdGO4wjqDEUV4eZ
5iOlILnvxBZ/vTLqkYGC0TwnGJVmSZ12ZMMQH3zxkXJL8Kz1JsugJbfQjSWslcFeXJ0axAGWyKAt
Dpspq2MjzF8xPqAdSMAb77oOS3fjEDxY/RLRZqdMC4DsZqS2vC3vIzoPzIYp2AlEZvZIOlUHoYkf
h2pc1e7z9A6aHHwBrDh76nTOG4p47k2JfgQ+nk87ytD0LaPpfbIo1SF77TPvBr4gyPMPQ9GDEO0s
Cp5EMUO+s+daK0CqANWFxfXVbbxe2njRtKczI/KAcvBIq3N40QUsJjKozx9WGBtpD7lzk41PW4YH
nRbRr8r9FgeLD9g0gHl9qQFyVl9H50ZdMnE7+jGEx07rUkj8wC08O+z5hphJvWqyhOf5PC6LieVP
hOY0tdyWCmjYZr0oagJZqfL2zp44FY1wLngH6Q2k1r/9Pr2jUwPKq+9twtUSVLIcrTLxI0Kskgiw
Y6A+QHtL0SuvlhQbfZkvIB4mf5+/KVzjpzxgx5gpWlDEcogc9pAfrikrr/rnjrOZmb6P5TUvIFDN
KYXEQvO4oYdhXLWmYrrxMx7hvfiD5NNcG1y05vaAZt2F+wSmoVpuNj0VFSUB0ptSfCaKqnNDG7+/
2AUmEj3mIjzDVoGOsOtHJiH9H5EOutjypZ/QV9wzpKBaSQf0UD1paZajQ4H2wrGZbaXlG8rOgCVY
IGs/Xu6IfDBCYmGdF2wRfHWshG4O34Ram73LFsA/zxTWv2GtFRUzjUUJYRpTn3gte4sLpkLEWhJ2
wgbkSWOZoNtuAP+kHH2fo8b/a7mY+ULjFUXJvXVwdew5EmdFDyu1Tq0Y3LHDiRrbyzyOnn2tePww
hoDrvRsKTvf1A6w00XYY7D6TrdzXPeNdpT2TRaZqz2gDPDgpGwHp3KPIe++KR0z4vhdKrGzfztrg
F7gRDztaEExoN3J4lci//hCLdufipyR0uUqdXcwMxmt66hOIJ2Mbz+Ar+JdV5BdhKDH0D5Sfnh4q
vZ8XVgIS7dug7/sWxKLnoiVE+PkZIMFJOvEMb5ryJWJJmCpBscAvpp9NrMeA4nYr7tcnlNkr/t1f
nqBaRN22UIttWFSuhhyFqp2pkXYXIEHt4/M7a/2YjFsEQuSbYfQcE5gV+jua6Gtz7p8WZpOsFI1G
SWUpcZGSnWpH7a3ReSkkwQpnT2CmVqYhJSTIgMowqESroBQwun7yqIMbDTJcuyzHUmvZGqQZpZRz
JJAZ+r0qjrVImji9crBJ4eRm80Oqy6XEBsJ26VK3uX8cNWDN1q17FL2Sh94GqS36E/h5UOQMbyUN
t0q2qNmVHNGkdqVMScjCBGeRoW696wruEVzFzXWc27L9YJvo2Uuoaja7rKi9O2DNDapCyV6TWEG4
3UuudTFYk2SghVZ6nZtUM6uSoyY7lAq5eE2QI14dPIn+O01Y5je4gZ5TVHhWqDsen/YA6BDIaun1
5SFRO/Al95mTuG8ejn6ViJkjx22hfZd5X8ovc+hhbTO78P7IEf3CswbWefUHkRcC/uCiW/ZX+OwS
Q45k8dMeZZpOFr0W6WWvrIIqGZsfKQ6XgbxunVW7nWMqG/AgBClXCO15mCI23qKBb1JZmcO1tOr9
77fv3a4rbvw3gZQe5q2mf73RQjHa/dIM7gboMz3AsjuMXMBQhlPfORLJjjhlZSb0vmqjv03/cZry
b0YL5DZSMOoTthoXZaJHnCvg5RvyVsyupk982YQmfimfJ6hu/fSkZ7gIlbvJedteSHyx7P4IaKs4
l+4L2t5ZeOxaiVBbEVQgZX8tIZ/20l+qwxDkoRkOGPoL0YcCsFRzYNDKj71erK/IzNU1htQuO2Yd
Mdoe3Ke7kBAPrScxnyM4fTAkuaNjWjaI+XrCVg/3Z7iL2slkBtuscTAhfuB2Vg3RtrJaoAL7kw/l
QACn0CMGBBrfAnyfPWem69gLUQD1OD/x/SputGoPAtSK7waBXeTF8Bm6SEa/XKTGk5mtw2QxofDR
eO9ynHmYbAEoWz6zBvE2ynpRU8floNetLSBvnBTAWEHBJAeJA+Xqby93H8+OxXul3UfF7vxmhr6E
mHzO2lC9sXj5Jwfv1CGf50y/YywdhfeoAHcvO4hy8cZgdBqQ0nwHI7ymbGCSJWMXqsa8rR9wmwtP
4dU9WrBpSdVkusYv3Gi/vyPZTdAQTAy9EsffYdnkv26QEcLaU1Xlr67AXFayKgcUBPgFEAqLjvp/
mw1kZgnkI4vN5UD+Qbtpaqr0hl+/bYZPHEPFSbcn+WRqKrOqQipWzkYQIWFDp7JVI0a24gw6gKqV
Z25PE/TrANtBPXzRI9ijTquNzojWG32rWF17uDbWHtFwHOtHnrqsfVci6sacfQzwpg2UkPzare/o
ta7ybjmFotE74xhKAqbSg6Sh3Kh5wbccZ1AqPe5pvB0V0qjo+C7ALa3EPnibzSJmMmMyR3yIMUdl
Cvk1E9p8VFxOkxBVb2LagWvO4TiqLrEFqmMfXq8zSp/zoNrzYDlx/K1zv9707gMez3Dbx7+xycZ4
XoD87S5Tddetm+J7fwsPET6wYdKLK9ncgSDGEKFzxEQ8EvvHOmJkpbOcm9atkSMp/HY63BFQLWUJ
2L//2ox5wFDs+be9PX79E1GUtK68H72/zXvJw6WutCeuqCQQTDNC5GrAeTFrKK7+PkDanUzzcZmP
WrROakGjClmU45TrFff4nmgGrsmI/ymATuFs65r21+TDaBwyYOt2iotjdWj3F5wn8r00UDaNQGD4
Sgv6F4g1udVRfSqklY+OQbhTq75uM8H25jxwO7cZubgyKKJc3wXfRtt1QqjuJL1Tu5/AqDCaD0xi
Wcs5wchYvDS5kcr9d1JOqBDJ+l24OrawZlc3Veg/rA9xZPhwYYQTXP7gtjpyJpIW9bklHoezWJAQ
/Q7iN3ARXo77XQvDaJfR97riXN1nabTbmOoGPklXbz17LrcwBZy+YiGeaQef7g0DmJRjytzBXjYm
OqneTTwc+ceplkwrY9JPiX1R8ia4pILOpZMVR7JFiuoWK+3mFikLGyRLTv9EpemKRZ1bC1TuKPEH
Lyp25zvWXuIKFmCRzztZJbPS3sk3hdM6aaLkWbZbzKua/BMHh1RAnLOYlNcxIUd3HJV0ANhyv3dx
GoOdv7XOyWQ2t0E8Ls1SoNaV1QGIUSX7dSYHnTCpCQVsb81dP8iLaVXF1z3lVgWDJcb6NYAEb4xt
QiW6WLSFM8iLqELBxB1OiJ3hVwkRRK3f+IJ0o77/oN6r/NSvPQAkU31n0+6mycqK9uW1kOQXl69b
OTRqyIIeTqSzsz3+83Zjbc5NJLPuS/9PqmcL1TYXMf6TdA/qKksLDIG5DdZbN2NmCGtq8wgEsIq3
sYbeV+MtORQfo+zudHUryy/ZTOgPxyPfK+Eqqz20Efa/vC2cosNyOEpn1EHPiHu1FrIxvmkayuiT
mJmkM6Sbeod2YgXiocz5E0jp7wME54nASpi0OPDLWbADr3OHkWjv/Otyzg8m2m7WuOOeZacDm0rZ
tGaZqT1Ze3bHkdb1VpppMB706OMeMUkPRUrnALwJl0inKgxGBunW9UrLouaz6X7rZl+x8XqIXggj
6e6uzsaWPILKv7ulmmwYBirC3PEZm2PIGSisRMW4I1aWa8lAu7n8jGfUgQ4TtQnwVZs/R/DnWb4f
oJsIZIMHqrKQmgAjlodpuZS8n/GveJX/D/d7291TyfDuY5X4cHAqmquoHxfaFznbbFIETiOqHAQt
AAkJxR9GtojAEmSrV7qGviqf9Fl+hiiIiArHo0frxfCjnTX8Bu5qLc6JOfp34P0BQqme+cv2Cqk1
whe3hoI6WEIz4B+b18etF4vZX3lJsjBg4veVqX5B+pbrs1m3moVbQGXjePRCU1TIHgTurUrGtG0/
mgRFT43FL5TQoCCkJJ4hwYtKdL4dTPeD5zBLQfhRrYH0aGAB/0jZyC6gbg6TEG3cdkHMRt8m/any
KJ0X/NsQNI6PZ0Ho9paVdaQ3i38bYn092olLh43RywupqdA1gYgfnjsiuVwiW4Ro9DYCDH4RzBGn
IrHRhYP9JF/ha7t+UNZNcY4fGdCE0wVRFSZhJUeXMn/rz2oNP1zhDl5Llyd8GkANmMIcfOGWDv1z
lf2YUiQDOhImQJ/SZlAg3dx0nwQNyqMCqOcW6xWoXzfNkkpNI/dqoUbEdaf8pi35AWmwQ0ekJmQC
G/6+lBb8Q2ChFef/qiTY2U0opVaoRV5Vpcuwv+xk7BsPHI69awFfRKpx50ScfF+o43sXxB6jo5Qt
rYlr07Ws3bvhAejgorlOMEWNbKdhVmLl/wAfy9QIa8G4dLDAWKzZPuUlxG9UY7+TjLelSP1lkIhD
FLOP5rNh0TqogPD8FEyFdrc5jlZ/YAYpOlkMqc54ZqTguq+0ObKPKklz0Y4otY1ZMGSpEecDAIqo
4pEpTn9CD1ukCiyeQ9K0uLxZo4dRf3WZIjRvcc+ljtTXU6FdPBXzpauI+J5L+ehl7BX/vux+xXl2
QxloIZ9jiQC2V2HRmtI5OszVxGLV7/82qhA7gjESpItyM0cBklmttmdAVzWUlwNJ88Q7BRf1pRGh
Vt39xO0j2TN/m9ONoAXO9rbSoSGvOH3o1XRDhoYy5Bzlq2vklBJgK1aYca1khEfPFG0QB125Jac+
1/PC9eug8oWlTibP/jaovTOvzVUyeGLN6OFPf10O9Ly9g25Bp+rvZiecRjZs0zPDOP2FR2WCWuEi
KT3EZKzEwxcfI+vZeH+8smPiaVp0HbBhnH9mfMufcHBDC+eHVkLVGQUXF96dYy0JLq8zCgMbrb7B
U/P9gb/dXoDRB8VcSmHGoKC+eEeHc0Jdomow6rKUSiZ4riJp+D3Vuz59BizNyc6q1Q06F3Ldbyp4
3/y0/h7K1yueQc4AcVGXymE+7tS4TVKvSUnwUZ7RE1Y/tI38Ya+of69kHryb3qOgeezVP8SNt8wU
oHXZBG4xzGalGQ3P+vVvAdpPYdqbI9aAW30JZQA+PKEb+oaBtpsza7D9AnleKJodiZhj2ntuPkDU
W8zo5urV/afqRNyTwacBbXnYkO/51Y7KQJgz5FTdlHh2bfol+dLQhLaEF4TVlTjBTAdEVM4RkYhs
nXO/hqkK+0hr6AKUrYw749lHIcl8uXrl6Vd6sJvqflLNXafrdNlgBBsq+q7miCcGspiWY3650vhf
IlserwECmnMrr/w7B6W8NDQDnYcJlBrDk0YJs3cOmb8Vgc+8MujXTKmZk9Z2thaylcnaez9CATDX
NgTKWjh122ugT3ee6KA+X0Vmh4SawP0ZSoSjIVRn6wgXoma22KLiU1H6WLBmBNxz2wpPDJ6s8NAX
NziKiVVs5hwk1qnIrKH/glOW4uSF+u4j6AQhAGmW49lHAVjiuDoYiU12XVq1g9vA3gZyY+++vn2f
/Cw8P4uMk/IydGhsNRjFHHSvI6OLumQK7f6sLuz1igaBOTTJatX0QfXKuI61J9VKxoslW5z1IbSF
xa2LF1HYFb9gALjECNNCBxLDPrlIlbhQ79+uqk8WIgxUbyc58kHxNYrwngiDoa7Ssf/F4zeCwBhu
rH0ajwtOV7Tzd9mQ7L66mQLtjFTOmE1RioVZennJCrk+GBhxCsEY18DjDmeboOhsgaAOmekJjxtr
qdEaDe37jjM6HBtvfUX09DGOh++mGO0vyjvkWYnioGY0Jo6sUavH3pJt075QR+NtjTFyYWx8jmnM
qtB2LGOi2Q5AORX9SWHMmacF+nYgR8lZywErBNZfU11ZRz0FOZ/XsefUdVO2ByviiBFeGvGvcCBx
bk+Lx7DV5n3+LZmCkv/PDp4naJCHYC28M7SpJSNbBV1Mt3U4XRx7Uujn8GKzBjkghDEdB3z5UURv
KOpCHvkXB5aQUYQ8K5mtp0+tzJ/0uup1EYk/1/JTgStd1rw+nrImPgs5vlrDJiMelH0Wj1+3G2zq
1s+wfs0in9C4R6TqTnPjEeIdJbWsr3Gg0oB1xWEr4gBlTGH56wqIR2K++JjmvZtr+NTnvb+8A86d
3CgLAqII1BylQm5gUSV0zE7X0lD0OkSJcsaVbaC80mR9bQRFVbXwFpocj5a5i327yUogOXG0IbP5
v+9cpUJ1MiNy1OX4DD6Mbp2xh9c1O7uE2bRCt6hydaQ7ooXrSlP3XRh3vb74juZi2MeC5Mkj3mLx
Fs4GfFW67QlAPwn1WoYzzdOn1r1a21oDkU6PhmDIFwW4IvyuUsqgLqt4QGBqgI9eToYY5gM8YVvm
y1waZgchnDlRVhyWbfGlwrIHIAEsgJRM88GBQMXW6L4mFMhK9TjXr8NM+ITKVO+IRAq1v+6if7Se
ljbNreJM36UYUe7FzRKUMuNGHorhR3jB1EvBgxxbavohT/tVhojlwhX/aTIPYcW6NoZVobUWhvwI
3r1lUtKnB69XNEg0EVNnAH/UCN77cyK2z70FvkYsktYIwBTwLl5Si2h0sjp3dgSodWv58pwNnQbd
sNQZLJPjiAIVjVg9dj61lp+qBcMHq5KooatfmLbOdP4lXqT5bzoHcfhaHIm+7Zzo2CCs9W3bdVut
FL7dvh50IqGl7mKUXNuSW53FADM5LjPeXhg35a0ofCr9O+dYL3C2HRTPKTkqmIwIZlGSMO/Mbebw
hYB9QxarxVGKWKOsUY1GUX8FyR9rvPDj86GbNU3uEXGopQI00TBuGSDnExaIWSkISUgRbVySMbeO
KPhCEa6+rzbhq6hlkWb5aKliJS5AAHJFrw/MseICwwqZMyUdW8LMIwkAIQX9WThc+DHmw75u2v4c
ocDN2kN9PckP1/qfZMjIHqM52hV40aHjSaCQ1BnrrDc/FKljqE0bEbVHn8M102HH36lH6vLAafGP
12Yz3/moEdCXK5oCn3nLF+rUztbP2llqIw04EB6iwaeA4QdsdfJVE0S9xcCP3ZM5dfGmJYlDRrXb
SwVnRDyKYu3Hcq/wB9Arhp/sHs+0Y0EtBw4MAKO9PLD//co3H2EkniuMiB3s6PPA4sMwVWY76Zhr
Q8pVBQ1tHoMetkSbuGKHzqMTsQ7/9F+lWRoZ8eOWh8gt0kMachjnCOsLQdxoNYWAEKtDa50bcd5O
dIZYlzb4rmWrlRJI6HueGeoKJKLtQrrQR0vtFFJttPV1/br9/F73LIaaeClw/gGRkzxmXK033BHS
ft7HVylqXfq/O3Yph4bpl+3FuozNtZjpTzGj1Q/hvbTz0JrCO6SxeH1cLtXdW5HmELuWp7I+Ka46
63x0CJCj6lkPr0oaqhBqSlQbpBB1LGcLdpMwBl0JaPajb/wwQxYRvb6YCnjaz/f2xXlOJJ45YztP
su62+YV9rWfMLhS7+X60couoIrDtAfZXeiOIL2/Y03u8C/4NAOk5AN/cZzD+8FRJTU5X83eDgrVz
HDcTeK8klcOynKu6Dc03WUKUp1MMEl/WCq1sf1aiTazMS5+lHTwVBJNxM/bdOFh9xDG2U9902ara
FdHKF6pXaLNHOA8I0YFa0BStalKR5x0GcPAuyeEFMGkW1lj7QpRLQv/TJhqTTpn0qKYeSWcZNmzh
xhefCoargeHsE5+LwPb2e3jV1WEgm06HQeZxlyKonqKzSPIjQmTUTd+jSco6zx3sDr/Ey7m9WeQc
Bfrvjd57cLH+pEclzO7Bkh8PVCZyX3UB8lnu3Ha71Bt1CLBsw2H0Rk8Qk1+tELpfX4kRvqXzXSwC
kengRsNi6fZyJ/mGwwYT8UPX5gzMs5J8DSoGgDWjyEPmNeyFU3x137KdhzskayHRNOTeOlAh75x/
46FWWvQu0SNoSCBu+onRpDzP4R6gKsYJrmkOSUSlKdykh/tOPlnmfMjyZjpYTs82KdgjvNaR7In7
BhQh7Ogg94xIAm84r2Nit5TOwSd/baAqQ+QaWne/2sv0C6QUE2yipgTz2SH2VqU2IirAI2RnM5nf
JRMbZ2gdVem4C0G0Qov1y7U74gLkdH07lBiV9W27+m4jluF1fVYBq7RJwIN5pu0AYEqwnbbuBgsE
RfmjjQmLeLlzQPoamde04nJn2eFccsDUojJjo1xdr/Srvv4+ht8UaIljNRDlEmcVDD6eEwZqe1Id
kt9Gh2+APdQtBm2LynV8DY+GjUPVKy/f3aP6NodbVaeXuiwymW5nkU+4/4BAG40Tdp8Abafo8o9J
K4aL79S9Hv9sek/hAjRJDwauqEVxmCl/+ieO4zJDFKNW9BDicpfMr3ATo8AgfWIAFo213XbGX+FR
WG8CNblhYuxGAricWpF5xCaYHKGQNM3u8AOzC3AtGFzoXtm8A0Gvgs9tLKBkrMVhX6LsWnIE+uQb
DeGg+9w7VgJmuT0o0Ex/5AyzU3t+UZNQrDQvFeAQGGSzyB0JJxyHBRWOuM6acvp+pLM4iwSWW44j
uJ5Pg3SIgHN0oiiCa4qrAtfFvRYMrO5+/lLP+ryAd8oDoGSLJtFL6TNJ+Htj71v9Msxtq0GHZW+M
Mj9Gvbs/uPTZsbEHdKkS5jrOzAUrd688NatKdAQxXKWy0iTotFvVTkJ9DxR+mAdVs8Dd6qIfK9MZ
/V37lxMw6igYnj4euhJaAKrAZSrhhoCdLO/ltpUBs7ql7PEuzp+nJy5Y52R5pXeQYU7xgLdL71pb
ptL6zpEEAtUn8xS//ByutLEdr6srQN9mL63Zaou8F4a8hXhIUiZP9sJCw4zRM8WQOr0JS2zpqAAc
WwZ0CPp5ESQGdwc2iAad55coiA60XQXSsxoKAta0LJQaQwpfK2OQ+Re+OFsFqcNy0BYZOe86k+cg
ikdu0NPlgsuU+GOaiPiDvbotl0+3MvafYFoqoWQ6VTB3ZooQveDV+Cw9Yd6dB8JrJW7zHCuV2+56
Mw7TCQDUzGhdq0q9OuxTDEQCxpQsOjZqtjWL/5UU3OFIQXSGVNHhrQ7xV4G0kpYz5UxqeESRHXfK
7gx6FPMGR4BWzL7Dvqm0m1EkPE4q+JoXNloXaAdCMk854CQ7x4vu5cQpoRrs9hKLySvlEbsKtPkJ
R8HLt2GNtFDl2KczuuHRlUuoyiSvnWHpBhR/Cndj7CFcPgSTBBcfFSrap9Zm5h/F/79eKQimpLfg
D2w7NRLLOPDvNwKG8TUYULJF9UPtLlPSPWbd2BRxnfYJI/1bRTvPzAiQd4pxxYs25U4b7osXnP+P
yoJCJGMIDmDbkyNR+CMGP54WfQL0etu9vGqXAN5592nNH4ILN6lQ4T/sT4RyOngw672diMWf1hkI
T5llqIgqAvNSn6MgrRBR2IG78CcWAJHkugXCU73quz/4XCwD3OPrRgnDBsNfacgj97AMz0QKh9fv
4yLny8V9yVXl3dglDXqZxpc07piTMasYzPS8OeD7WV7iqAqnKCIg11ryLqgzKDpELRPNMotycjiN
x08NHf8pXLpJ0XK1mIA4sMx5/L2K5ZFzL4JbMQ/0Xw0DT6tT2LiWAjcSr3TCoXTmCDGqBlu5vFWo
2Uw4sdppeAsxvgMQpALTFnu8rQtw6RRhprtUrioV+hucO19t775mZ/9qKJLPpZfN+pvlGsBGy0gU
eY3xuufHvnl7L0Hm69fm8Kqy1Ns6XjD/v6P1XPBMC4Z0+AMVS+DHrj+NzEDh5VYfIKM1q3wTTz5i
DCBYHd+bGq7ItOcZX79BrTIzh5xaiiZacesrHUO73d0NXRHONapyVVC4S6ytreUbokz1NKQFHRvj
8MN9bDsuf2EzMZeCruuQJ9vkDq4I2EP4TqayOd9Orb26BpQ9t0zcliXnPYN/JiuvzGeFjGiFZjLH
JauYSRoMaAcezsYOErljgHpveCrTRfoyjhLyXHf+jNPYg3a6g+z/iuLJaFRQiYiKJs3GjJq+Hxw1
HTfsXF3kXmvHYEuvpQt4BaBY3HcnvHA03rs7Ryv+MN23Zkef5thFpUJUkD7yryG2Mh/rO0RLFBpY
vLE8ZdHXTTnghmPcKulBa5NC53bO4MSOQTZGszlFwIDA7quhLcnFOz8OmoEkAY6M0FGtyvYidj6H
u400ldY1t4vSILGMSmGz7CC6QGhawyux1mq2WZIsh3KsnLUzSreL0sP7tXy2IA43NZmNYhbK2PZA
8s8oXT1BDeRkH7EHZky5y1sHzItNzTLsJpzPt+anyumoEFIXwN0sTiGSC0+7AeAE4j8usPmdXiI4
9OJ2RgxR0ziHM9ADtWj78aK+yQFU0EINcDvwbSO979SNvO1p+Wbvh1dKTewx+lCPOlhEaxCpBfqs
DxGWFi/KGC1zoDvdlAvSHNlCtqgDMiRsvuZcMJ+nk1QUex2JBwY7eBAPLBBCB0MCG29kMtD4RxSP
Cym00nhdw/0T9qRGb9UDukoAXy+UUJA7bPY/yZOgPElZ+O2O/VsMIxg5HysZO7jXwT+mwLd2UlDS
MWYCgzmi/0QKodMzvjfclV5fuN/14L3CIa8Y1fKTLnzKADSs20QrlCC8ga172V7YQB0OxcCWJe97
K1lYQoYlmeiPhWtkiYKSMEWEQwW33N9Eof8vENZk84jPBnzgDXYtNcgjpCt8P0bpRTf5PEih+Vva
986kmeDTAx2ioowCTEklvvPo3Cxls9xusdZVamYkKiymfiG95CIZ5CsuDv+Hlr1gDD4KYA+ovdIq
dLmf+mhYnf2wpp59nghHfofFfutlHtourx22tnh0G6RoCXa698YevkiN2LFeu2/2KzI43g0pw6bZ
OXSKJS2Y6eFFPJqJN+eUs14XQjMRZW00ZOVbYv+8MROoY3HCNDGRbGkFadcPyDwCvbQPQ2DFQvpx
WDekPZfjzEEJ+hEpRY5d6UXiie8f5xBwZ1RFP59MpevLPhsTSC/jj3jlaQvHS0Y3izd5gWG8kLis
H73N70wwek/ikHyJwDNDT5bJobLWVKitO3Rr2fsuJy+GPec0Fn9UUfqg240Plrnw/qnlr7VxKAhj
9JtDFD+xKPrwNLGGT4vjPVFWq2NDm6wEY9hGJLWvjN+OTjFNDtW2ViYsHsnzYKySPNKVVnKHejmj
KCK8ixY+W5dY+Za8+vvGIeI28OYAZ1Rhd/Q+J5wrHlyZHHf9eUubVBiexizPSzAJPgJYbfHJ+mFU
g9AnRmldBP5KhD/9jcOfvC/gkqCY9OzZBC9dq/XFYawuMeUin2G9dja/wqlW9boTInGYX53etKQN
iQBNS6/L6XIAxqCXUy1rHtDwBsXKAPkyMbg0b+1V7KQct1SaSXcmBLueu1TyQ2bEkWlkDeog3FAn
YMRwFiIMoaDoj2bonkOP7Ua14M2tKoMbLziKbImfa72+8/9iTWRdwbUkXOhb7D0q9RiHBOQ70yNt
dF1gRkB+F6SlJH7uRJ/cKDJ7uzF8t5+4mnB6oGK7dHxQmrcHA1ApUjCatGjVQkHXjT1DKCPTyUhe
C4KQH/+UdSz/22R66d7JrpBS90p3q0T/E9c6hWcYI0KoDP79Jz5lSa4xfiVPa6I8+QMc5RmKEFee
6ntqVdKmMq299OpstKHDYK1kSzUERUgZeHeeYVajg0oZPTzfPfbbBeNoOC5USARmyIjroz9o/RtY
WVa0JGEq+xuLtRbZdBPHmG8ItSRsunmPQGVBvoB/EgpzBUXFOG6yXuyk21OGGjiASaW50TUaBcB2
mxjy0ZmtFmDBx/CdxnmrGzQLJpol3zTVAWO+MpXQ5y+x5QHgAoJHKOXVYHp8qY3WmJhFZx46oJFT
n46HNwHrZpNtqN8C5Rk6FgcQ+s8Kc/1oi0o4PJzo0CnI7UZvzaLplQY6g3PTvtYmJw9yDvRvUsk4
gMAJQ0TnRTqkn9XXVK6Z0DAe7ZQnhowIdjUW7Fs3qHCVhQbNEKLtEhmw7EDgT3tchmvMYL2EJVFz
b+W3fTBUqOJ6nU6rsmX7F46hZsI2wM/JawydE+6lKnwZey7KnVQNyqXikK23S5yu6XNdbepUFopu
fK5GgcP9Gfm09+wKvxi08fT+tSwKPVbnL+j93ELO3z08NTyt+8YifywosKA5llPM8L55Ng6w0sDe
EW6s+6csUVcDdEFjsA4TfxZApJSa/3vTm2Sr7L5St/7gKvv3C8tvJghdM5fmF6ip1vENPWKNfJ+b
Wpihha9iPQs/CtxF5h3lOMvzUSKIZOzziircAxEhDeIwKUThoahwcdYB8241utB0oD4oUElPOm4w
EMQyuOsIHwHD2vG8JULgqIKsoBye8nwXls4BAgJC32UPHkgWkhmRNoCn5iIUpz3SPsC6Fv2TO8dM
wOEiWFKeF2+hdiDMlWLpeqFGCpBicDfPyuyak1h3eYY+2QM3fbIwf6U6TfglFFr+xHqQ0U3LFDya
CKvFIVdWewN6Mik3pH2/qvh9s59uYMFACCeP8qLNaJxrGp/wJBSezp6QIaQQVQ8AIGoSNVY/6ltP
2C/+qGYSKOVaEUhGC0jwEVHdFNh7opGasmzeK4dEjLZwzEhFdxIY6MmYJ3vKFkSIrwmf6n1N+eDR
SwZ8IATr4ohYb29R/WS37Sqala0bmeaPEO70LknGJSRR0LyunMoH1GVNXWM4DCqkiRgj59kmr+RE
goz7mAKT+YzbHRk9AHchTnp0mb7N87qea8pwGuojZAI5mmknvwNPzo5WXSe47Kge1GdyCf/L5l7m
kSroP7uF+iZiF4VFGk3n2forTdIf7sEN6GDFMNIOUzrpng1ss3cKu9YFAIgeduDPAQ1Z/nv7ZGaI
ENKpfAFwJJx381nLvyGUaSZMm0ogliXnTCecKHtD8l7n4MC1EquD5n/LMJqasgvrGOXcl7lfCcoA
qCztUxPfpYktqtrwEWmI/cTRp9ZxvIxI8EWfucTqYOnQdrNgCl5yfooSKO4lgmE1BHCjcwXHp6li
/ubwa+MvhuM0mlgVz9mnSzDJG7ZGeIDGvlTDMdIagoEmc1PMTAhLwjFZ7deibQYS+Desnvg2SqI5
zyj/z8jQxREZLu6MZrpz5dzLlEP5cwoqHTqpuGkK2/34pUCKQ29aWkFCxyTASizOZBecx6dlzZEs
NahtXeOk8yqgXOgm3xtRkNUtV2iw1gaaV32L4IPV9IWYDbyyPvd+oFnlNdzILVy52PwSn9d+YRwv
3PDMWBc+JUiSsTQTmATt1EXZssFuqJanTzLu8tgoHikjdb7g3ryl2ks0Dxk7uEm9u/5XG3cWiO27
4X1dcCxfiMRz2Y0aLv41uEFgn9iSQ4cFUUjpdm81griM6+e6g+S2D8Q/7Ev0wFdTD0IWZZU1jD2V
qelAJdlKcVMNIyAuyEbvly/3TSPGG1tqDH9k24qiaMi54gYvFxmGwpW9vAtuhpgFUt8bKRvg9/bf
JcnPa2mzuUA+V9OqzN43uGKnv8y0Ykpwmh9Sz6LnmsJMecNDfXG+iosuyspYFDrxFbahOQZZCStn
zji0eI3Bz/3frMBsARfkpfK4CZV0LVRYmNyKOsNFxFR6K+/AdJcvB3FqQsNKdTr0l/5PUKEn6oH8
lkY9I0L8JWLCTREATOO7nS8XKoB1Ad/bxhACeVHbdKiJaQPkqDmhUlXsZdmn2G48JKKyCsD4L3DP
n5QjVom6YDn/bFJfwP+wGB/VXM3BQ4gwK4Q6cqlNzSHvpmBEYYuk86OvxKg8EV1OvTcKQEOu/Aep
dOBVD28Tpu2BXflTe1ZxUvwLymXOv10mt0fZE2g5tcF/HVjBfJCGc04h9nPH61AFaSPcVDqUv+pH
cSrLkOpSmhFupd140n6Q++HMO8Hq/Ae9TIChsSMb9u1gLpveIovnApf8Ll6HuZoGOlGikPS5P+Qm
Iug+Qupjx+qUodXQ7ukoUPI2RHFbCR3JUquseI4C/L5OFQC+0FCfPRKY/HpJZN2AqNnhEXnlVetn
9O9YEbAiPhNbA8wGtLLAM7KQnMPoSYgRI0oZFXgCkn9gDnh/4c8AnjUkFLiYkK5OotfwSJqWRC7g
LTq4+xESR4s8ygj3+20wDCPsu9iIwsIWKzDL/KGc5av7K/n0F5X2dE1spkCmRlkBXNfxOdU4XtYs
G617iLrfIQRU5Z1c9BJ2ZWHu21wa2PExO/czWJ7QRrGfe3V3y4uPDvevglNRO3mv+6Sf9I8NOahb
XLOAYw4obK0B7hasFstAJ1aPhIjIFCZC2HTtZ2amle6M2yZktivk/Kazjf7PP0FzOZUWVmUJkubs
AVEOQp0yJ3Ee2ZajjOfFItddq1epF9H+nMZ0x7YYCPZ1IVbwZuIZBwPW8LgpdVRRciCx6QNj2mRe
1fnzxQa6MN+GWLfcLeCbHnO2ZeVXHSgGMqB4T139ChCA5Q6zXEKY8tn9GLw7PQSZWpsPxny0DCQW
4UScALR8EjDeUgb6Q+zaAcSoC2mvWmH79J1d9mjUucRUyxDE8wiNaE8NztIgThOIHh/nINzBK7/P
mU+Z74wxUnJfixjQL2DL5Al04Wla2todF6me+d4YyhwVTlhmyEoagsJRP+M2SeiCpPWdpn0zNEUX
6dsso88nEOJLbEXqcW3WtNNt9anl5C2r+JeOYkmQXuGvLE1yiOyBMAvgILBuOVi2HzUYyRniJXPM
PdmkaTMEtCPe7yhNJIsolp29IXYOd+K2jUCHWtwX9TMwSxGZAtyWQ6FWq2yoJf1UOG1sbhKeRpWi
ikuk5G08Udr+skFNZoBEQLRiD0639M6w/+KDwDj1B0KXa1yPwipQHAmRIDqXQxAwl6AQ7q24dZNt
9PYbg+x3ClfB3dYrN2oqB8XHhJA6ChTpNQ5rqlJvW3Jr1EDx7j//COQdXuied4zCbBWO1ztTfGJo
HJ3oiHDfxvq7oP5IOSG1MoEL2MUGxZd/TTBnBulHks+7lX2LwiN67jZLXJPZqKX6hklds1S9q2aT
Yovmil3Y29C3FS+t4h/9SYhQTs3M2p3sQzvLSqMbMnPCzXECQ+OoeN/dAtE+NNLsM/WudNqDzffg
s0r4vL/TExhy9YuBNlUhi4+leoMZUKK4BjBqFGF/BdVmRDs1p3PZcIPX88qqGBq4WAoUfx6kuUyU
6Z1MfgDMIm+KwtiH3TedC/9cxowxY0spG3rYz5HqJ5qX4bhrvH8enB3+xALIv4tNJzbUSnwMOFL/
GMrgbHqVBMLtc6cWFJY9mtvq7rRhlXJiYNe8L3pCnaQFkk5y86+oDlrtef6ilgk9L8veSMXdLVuG
yy7DHmMKpzJ7BW728plWM7ac+o6xp/Sum9QueZy4yqVCi/1mu2glhxrizNbrUd4wsZnz/s2Hfbtk
RTKVANLsgIjK9ufU3ceIzXnuzBY5OLSH1v83oJiXu1+maeHKp7+48FqUUtPwhRj5g6O5KYVxJQS3
GU8f4ncDl1NW9ekWirKm43gWqZu9NxWwaNG1BZaEMCLU6Ara5DDSXrIV3gj2FZKPlLi53x/bE+xr
f3xgHLHh7AE/y3zy5No/5GKmBID8bsSTFVaNqKbiGICDDBUlAvRlNLrBJ6zoNqW9RNa2kVH5Y0Mf
rAMQ7K70kKujmTDMpy0/thskn7+g6+/GAAtIowvBzcfvJD51orWzovShcm074jfZk9Zgu1k+FUtf
4nXcAtd9OpFaiiRu+oZ0i3yug7/YamuxedES8R/NA/z+oO8a9RCfR/st8xvA3LPpZQUdOnbN4EH/
uwNe/6l5DAwoystUGesrS07RjcAiHxm1p/L6xUN4XgnmaZX1huZl6YbI0vmPEgdPHQ90p19ahQMC
kCRcSjHSUPEVXbJrnVIGKNzVS75+5fdofhjntkjShr8omdp2+SZJfkB8mmeAamaLN2lStjCn8r6q
lGMqMudGJY4QicRTAm5GUvyW5n095VB/oa2ZAK11OG19DNehCVshR6eIdKU7RtQBgfiDMDtv1Pa5
o0yL0Elp8cR5En2RACLqWJ3Hd2kMVPWxSjuy0WJscjzYz8g7v1sttVMX622zWjJnWIy3dZA2UByQ
OkryUAGr6x2ydrT87hfkC308u8TRiQrKoR4ofeCymQMJ46XwTAruRw1yxVshQdluTgtIvqgTYk+o
YHpOyFZjWwfQEbN1IE6xrhn+593qOR1lN3hZY1jSV0NNM8zjW4AcWA+JQ5qj1ul2R8EA9ZgUdEgz
QITZRXN1Kk318zQQ3HvX0fXh0E+iVA15JuVU9ScsUphfjAfLlQ1xjWH4H9eMhtKsvEKitavPir4M
CKocwu8OUnZcEmPe9IKcW5vbuqdJODVCp7Pfr7682TWQ8UcIFA7n1WX3R9x5LU0h6p2xJfMjPGlr
1c1g03rzzzOEKgS4pQsimRatWfKRonlXIxsTW/0ilY9XraB/xEPZZ8gtwRZ+lQSDblsz1xNowIwA
pVxHIdRtUFrC0CDIZT/d8gmJDoIPw7NlomCd1Z+1U8aEIhYAVR2JrutUhwLx8E8bFu6oDzATrRF7
ox85GcOFlaEEo2nfGAt7lWs1PT59QACIGOXvHrNUWSChQsHX0gBIDDZ0sAXNraaeAOunzsPy2sQ7
FGvhKl1iyGmEL6rse48vqgda9irBQxNnlK5XUjiqyU6FOXUTgfFbkd4Q+Fyvo9T9boaLQMIYKupN
9CQzD+YVSxryMCIhtHYftA0zmaH4MS2bKFN6Xv6/snEAj12JL1WGqMJsn0vxHTlpLMu3iV7Pa4Uz
0P+rY77ylTkY2AsYqAw6ZNUlXjWSYBtxGNy/EWwrYecWn3Ez/xPEqfP4QLn7LFSYUmLeu37FMzCh
QYiBhJilJLYWqyp/F1xkEc6g/ePqUoy8Ps59uDmUGH54zUzqVcmHDjxzHD9g9HHXeAD3aU2Uiw4n
dMQFrsAnweCi8ZwYUq/wxgSiS4FPk0wbuJwht+QY1IfgKcs017IAAtMM9HcVf0+tsRMLPMCMqOJv
ObP7kLiMfNcel04fKmWoCpw1dIIssDQk/T/pEryYUOJXfwr/naRCO8FLEAlBwBP5tlvcxxXJIv9Y
m6Bz+l9flVzRGsB4nOv+ZDRVkaeKtGANj2J2znCjQ1ttFM8uPY/LqeWSAln66WYFu5n9sNl50kdt
jrXNfcNBIT/QqBubDaiQkJpHYmX57GIr4yuEyFN0GklQKlKyfyU9GNXyPT1FwvBQ1GIW6LOvL5E/
+m72zSsxGfkLy3QhSrRPIqToQrZQvRods3QXnb/qCaboCX4BD8Kz7KQm5pmoOA/kW8UTBN5P31kN
RrMysG1N3GSOvCkwYK1N5nUNQ7ggQqArDDlR3onTAfOhGUqDqYeSXjmQptIych8GfZCjrbZrLbyH
SG6N9SMrIv4WqJ6UxHMDsnLBTXic3cmGjd5zS7wINYYafnZZCQTYrzZwAayaNUOtXUyYxuGz8er4
mvbX8NQPdCkxopFq4ZFtvcGftHBL7OJ/KbIsf5ju/JArnpu9tcXCO8Ppa8NmE21yH6BmuKbD0m5U
axsdRiMtHanOBg5SJVbzINeWe93NPWJac5rJP72oAvqzGweT5toFZkQERZA0YuWWyvC0XBnW6O5W
8x2Fbf2uhvi1hasY6Aa/80tt6uTn+0BhH6Grj2z0Sly6W34VukxulfrMZ8mPQiGo8E8NSfH6L82e
FS+s5AtJoF3kT4nOv/rZct7gE7RRrHJpUORxoIaTB4RWhpLdMihJzmQLs2vroi8sH/GIIbYPsvLx
4XF5T7uG3Vlcb2JGmz1gy2C6jj7lVKdIjk1+A2GfqiLxrFkGsJJ4ahg6A92nihtFt41t6ZeQiKUW
wdrMDIeawqjkrUra4LdUjSvHX97wJD4VHMoRmhcFQgpXyO2OqAVwfiVTnb8WU6AcP18HSf40ctDL
qR8G0UwfMbezS5xDZCBSWRy6XhuRH77DR1SFDLBPfM3MBM5DJPA/VWxZJR+Z34zOQ7tGz6gL4Txm
sl4SJf3BQeLbiKJgx8rMPRlUqsYxCo0EV8vzhNYK65x78LP0yBks2VePgxb9+ETuVj1m89iaOjFJ
/Wx7luoLoT/sdC2ZReiuphDW+vBMFkovyxHffDRHKI3sH1ErSy5fjGhbA0d18UbHT+EXevwSjKKX
FQ6X3OO6lHEhcmzC5uE1Lk1t28sW8OqMo01g2eFepVi3qeAEFZ2Pw04yqCFqIXUH/Bk08KnTuzLW
djXNWIyHkagRs3tuEqxP6QsjUqxOy0nwqEbIjFvXp0ocas3UBBCoHSOUxYAkgqCH0mug8/2imCkq
BQRw79qJrIT5QV4c1lDUdP11BEFbJVOCRyN17D7iNQSrcExwbckZ9ShXAmeRjHKQDZKZxtnEzrq6
27bubUM1Cf4vumhOxcS+vvbFUbYP64qW8dAxmbd+KyZ6lrRcPiL/5exnTMtcG9UmnWKyUkYh+IMh
0gF7/58J0biMbo1PAivnFg/TIfxdjJDY7VFb0kxVaWOsxGXY/WV/4N3LUkVu6kbL2OOB5MXvQlJ+
yUYt8HF7SNerPHYr6a712JuU56ac9h+gRaM/4ZWTRuFejWT0vTgYmtejxkjNjQoUOlIYN4QbyFM/
8s7FQOeqz1n/0Mrym86Pvg9aOPR8QwbBh8j2/b29uk6Mji4Og7Ggu5aSddHPXVVs/0fvVkNAD8W0
FWurDvoHO56R7QnyaGQpQ6ypvp419oPJXNmjaB7zly3PER4QUz1YdmZ6W8N7isnF2W0D+hA01mZd
wC/5878aFm2FDmKSknk7RA8rzR+HrHwmMaahEv07wZsZ+T3eW8Dt2sv2zaaFA2dfetAIgWyIEpqz
Q1W1fDjT+EHhr2SvCziOs8/ElIS4Aw9MYcsOgjM7RTvx0fL/oR1NaJyYOtTqf+/DrAXjN7se5l7Z
XZHletGPMlhCiSGDvLvL9VpPCfDk/nI1t5hsq/DgyJOiiMvplXY4+iO1hCqcKo0KHGfD4w5jWRao
PHHG0leaykyn7Mvk/2d03BVEVxqPB5bUfGbRnXJWDgWBXPCMY4PIoEr9SDAjnWCoN/aw4VKnYgN2
SXS7OBS8WZo35PyBZ6xn2t3mD/PwHsFlVlfLAQ545jvYJ4Z4sq9INeK6M8ujqffw5Gs84cxvORRn
vOZ4clxsLewccJLwkUUlY+ZvCijzSPhUQufFkVBgKt685iTNBGYDFUkcEZpOP29MnWLJ24Iy19Va
c15iRo0rCr0XOLDLaeygWKJ5RospYHltTm753/2QfOao5AmH1bUSyiER0CUhC2HKNovtyiTdmie3
lJt913kI3KZwx3/gtoBQMM382+er6ablV+qd5UnBUUPaknOcgIl6MAdbC4sFU2CalFcZK1uKuHc4
yyqO9aIPu0yUpbv5FB9LSGd1+PM7/sEVz5vzoPba+qQpaQ1+1QFnfYbOJ8BPNMotVgfyFkKACZAq
mSC2AzuXK5BLU9g25KU2I+G7ipbecSF2BNIwYU5Qe5SAyU6rmUbxJPYHfdMf3pU0AEED111fbnDa
LTio7dwN1CmvCRDEVfSxQSkbcdH9v0NtUfm5s4Cuxy2GDN4KTAGn+qozDsemBAd3DvMyMR92THOq
/nEpk7+/cII/e6i+NThkOFScXVzeR+5gyfCqaJoDITNlCz9bW8pZHZBnJFmN7jAKhMhNg4yIhrML
7EvQFFxa3ZT3mL6ft5j8dFhjAXj2A76hE1Ze+sbORg//QUMRyKUSIR4KVYp/GQ17oGwWBfgQrEdY
B+Z0CJgvtdEEWPeN0I1pYUmAAR2uj1UBQIDWtuGNHhRAGW/X+7mWk5LYqcfloMLgkiYKYaBg6O76
HpHBUEK1vl09XmhxSlYlBnbh2uigj2p74RlHVr+PphUsBbr9Fvxw+nikKMMPvIi4p0JmodAgNaBO
T7RREwrlwFI+NusMaBDSO1ah9BY7igrvzHCnHX0fivoC3KytbjXYwlGPKB/lr9UwiPhAezTDzrYR
L5qyuq/YyJvoNFEA00wKlfK3ole48AxX/YchLRPOR9p3N1iIJiyMFKm7ua27+Cjx/uQxrtLMB7/k
YD+Lc0NXSDDi5n0t4xYVrJfdJujVSUS9qN8rJgmEt+weSUIG85HFgq8SoMmM5x9rMG7d7jaJ2qMs
kZrTzRfcikqHJHElvj7A6IAWcOD3maJ7D+41g1WUdRvbFjs1EBv08/r3eDXBSCAQD6SU77E0gc8L
6jHKrwtOIf9jC3P7qQnRAJ7RiMq/8Bl00KzkaOCdpgbuYU51POL9h6irR2FvoP3alR5/iJBeYBfr
/t0GtPjc9M/TURGjMjX6b+klauZLoR6YSBXxs+5+UhxOf+tJn/OSmN1grPAUB2UYUujT7NoalRRd
eq7EXnbUC8CRbeG8C14LKjeuimZ9d9lzGlic8zoooMfc1upYZ7DLfyrlAJ1pidPShqAqWeot4j65
PY6NokAns8dnu2hl6YOkuew9SGaIDYM3ysxoc5XY+Emito3zSM0Nq6dqRIYJUlKQN5xWf0aNLIpt
X0Mn2cYV0gdA0VWT4ut+HmiqaXCaT2p3tkNGs5hzAtjHIoEcfoO+6v/j2ala1oj0kV6kb25eu+Li
u0XvZZmaxCWI0VgnoaMT7rTOXn1hRuPN4TmnXF6GxQC3TmPgafqWsJRz+u4qqUldxrwtcq9++YCo
pYCw0ZppOP/NhbRFpwxhsJFVwusmG0YRfMjZy+RI7x4OUL7Thm2hJmfIwhb/xHPxNZNBJ5Zg+0g4
utLuVEEFVADFrTNLHa//YNkqL1IHqlZPaY1Oh6H/d30MNFvBOk/10rCNeqbUt7kHgy56nQmJ/LIB
QCJ+87lHzC1ni9GtxVBsz1//GxgY7wNcV00n2JipqnoBtHvV55kb4kJ11HHfWe9Zxo720lcP9pr2
jofROuCVxHysP8RzQOwNK+pJNmXhlhS7L036763G7K5V6j7wdAKPgtFai2ueuY4DmB2scR79QnI6
oz2BOFTTZ467WWzxgPxGmFJyWLBdo5eLBqNyurVEzEwfg1neFKNtluutohjrQ/iiwcxzI3bG2p5R
chNNfH0tyE6baEZr02teXItLoMtPtt48msg6KOR/ZDf21uImZus3Di+f5301rwrZBguYtGivUOiU
0IPhqdSgkQ/b8v2X3diItGNRgQBWGmE3uYKcAQzgaiUGW3NLIHGiWG7nRnMp7/eB3GCyAR6IizpX
2wIyQ4QnPUI9no13lwg/5Nbxq2r0sy49asTGMhjzwNbWrtC/GenFIlMTVWUq68X60MaLC0HpH6oe
ZJZtf2b+QQm/6cjBlUspY1lssYQqk/kdz98XBP6LQcFLISX3g+w9gyOKBgukw7uxqdnjwlZhx1yI
g/eJmuasAwGiyLoDVXYhNM7brVMRlhntvq5F/F7d5ulrmC/3BvofvjHXGnqv7KE6masQy37Uq9S2
DOFYZoPfz5uj0ADi/o2jNb8mutiRTvPlWeIShDqAyQv5cdgVMMdJqWvHlpzja0MNE7zkatsXZ10N
+brrGp4dDC0e39bLj9QXvPh5X8D7FstmQgaEprCYMkfgGGCKD305o5D2QjEyW9p/S7V2e7l82osS
ToHXWCG4WAzt+bNdvBvWwsjNRuKZyLVKDN3XNvuop07wyPrwVIfGaCMov+lIjDxY9P8m1bHzHi6S
Z06yHkEre4QmJFgMrjNhoQ3zrVCTgtVVrWqnBM5G9ft/tE99yYe+N0hfKCt2+6AoS0Pz41joDp4+
A/EzAfoaYxLTmc/AgU2eb5yD76m0S/tvAAChpC5ND47jPf81NU7MWTkymOIRGtESgjGZmO4jkdvp
3IbSQ0wl4pwzJzhwJ1U/15J/SooEYWVMEzhu0pueK51EmIeV7+8thM4nAjwZ6+q5YzVdisjlbcH+
0X6YJAuYSDxGw5P2SwgtFPCLSt5VYDoA69/HmzBrC68HgXrxl/PvGGCKy53AiLotI4UMCQrJjvtq
xyR7OPFITokzKD6DH3ki5343unKuMnMXY4CbI5ow1Ohflc1xo6X73Urfgx8gne9GswUEFeBtJh+P
Q642Wv0b0cd6bpSk77tAEpNpdIcpnpGg55DY+1DmvNAVAXzE1RKzNXmDYUMg4iEJz7vyb6T7wzkm
UGPGE7eITjTeJpX3CFNU0Z+lDLHSjsvTtN+n7wXQM7Rrzz8DW/6dDz8S2Gs3+EeeauzWHGiQT2Ix
NTDN0AjYuxGNy1SOoTwx01oEMox/ZI9S0liF6ytfIdyD4y5jP230Dt2oKg/DyJC2hD51r4478W9N
nQcKrw9fNlhqLUzc76xy/HEWEgxF4dxSseSTWL5z2XK67NYiPbRFfJDjJ1MbZ+XOLJrRhzeZNe9/
UEREOR08IImQ1/EV/R3EWO5qjXbnWgDrkbQUWGg19CANYHiJJFSmBhB47kkovY/BRXwCqWslawmS
i84kS73AsMJyXAmVWFQ3m0xWXoVkxzps8xs7vrwCFX5Zpo2TX7i2YxE/rk0T1MUUKpuEDqdLovnP
e1zOa5ODDtqrZEWqPVAEN9N8RCyHOL/lzVSGXqrhOf0tg7eH5rnxwIWaYvr/gLWsiIveO3/RWOEc
i4JzrN8vJRMsGxd4bxF9KUNCY6tAv37ke8qDesH/0lCqd7jqj7GozB6i/jVyN0NL1s+NNgX6jTjn
iB87WggPO7INXhmIkgmzoHXGqRIHIyTwoc5CfDIYLC8QTeThurMAl9xc0TFldU/eMRgS+qOju/7Q
3Em6+jMk3NW6aL79PA0mw0MQi3kgSNDKgaZiKKK8OZ0hMv4bM5YP9ssm6yYNEFdMXWMdqR4WdUCv
cS7pQ0d1ye1nzcUBTiiTfndSDP6v8QZ4heyWa6AHKczsJqkPKl+9wE7rjRE6JIAEz1DZpW9pFP3y
kuRZHUNFpEmhaMMzlWqyggDycANxksN7GkN1tsV9p6UmC6dK79NpkER7YPz2RsqBIU2asqD9yrwL
KWZThlvhqkvA0B2lYZMmeHY9fQSZ+nMjmNNimB8ktcW78b5EmCrYYw5BWiSyy0Xg5cBie4TWaodw
oNA+qcvfAjFFiAOz0xsK3SeuxHXulwRKUtw0LMGpBg7xi4BU6/uXfzQvNUsmWA94AxIlej6RKcOF
ZWhUcSae4Pd2D1GWjFP2+BLI9Z99N57HMBeaWvASFM0AVEDM82sVwxKjg2rKPOj9hCGKIrIOJL7Y
aOekuA5CiYACQoYiIQmrEI4EGVIa1Qx1GUldk8Ylz2hkJTdKUaOYJKg57prGstBTfWvYGw8hI8HO
PmOQ7St3BZL2WDBJCPuQ2yKYnmiun76TemeV5yAiQEdoXhnIPC46xJReKjKuxp9aurNrt+c8fdtK
nZs1jBca7SH45HdG98kJ7C8PgqT5MzqMpPPu1TB8FZM7tzWRCHH/fcjH4W6z27zLsMDAgactTFMP
kqEivJts265vkG/V0truuP80sVtNzym0R+W2V6z2JxczbFO1bEAVQni9Ji/Mu228cwBxJ+HvEnMz
ehaMQHaWOjD4BLbRZsgEAzR52ekB5Q98YK3P0ZZ/otVZ8ITkBN3mwP7ddIjYlikykr43OOpbrA26
a/uolVVY2JxykzJyzf3Xdh7oj9zVaULSgiR05R4QTxuyIcpwjvJKu5kDPZCV5jCI2rceAh8rgJqo
kDKB0s87FMxZlBGElOdkz4WJ+PZ37/vhMXiZ5wjh1GTMCKLcEcKT6tDv6e4Yz4ZcT6GkSjxB8EeX
UHuJwjGB4FVl686qRtwVPfKJZNIc5EVfuooH+e5pP2swow7MUfQD/Lb5jdVYjrtH5z/e0Xl9soyP
6S2JZfJd6gv0zVvZOGqJupMOM8PvpQjkfcexn+qUlDEYtWgjKgFZWWZMtfn1qbwGkha7ZoYHs3ks
clZMkxDZfFiR56APtPxBPGD+5v6uXzt57KdVIAcS6u3ilOSDCCSaKYe4P3fnHzgdLK+NEq/eROKX
5lBxiMLBHZlFBC9u8FMnG3nmctvMPk4+pW+dUy8QEEdqW/08Nydv6/oH2iKMikgMJ/Rk9PJ8rW2B
skGDtyhJpLfVxJ0XDewSLxOlAjPYHdjr1cJRuSG8VcQpDieKDw8x8RPjFhxYe3xiAJ79J31+iTZf
q0/cBsS9ls7mrW8zFrlp/QjOyeqbizcSG5jvAt7XEAqP0T32dkn+GqaO9VZXLO2Jz7mrVz48dLgm
ab0pauFQ1wndPguQqt0EG3zx0YyGWf3PrF1q9gt2nntDL4+W1I11qDrH4kozAfjl1uROjRbpgfB/
fv9WyKJGCCHXHIgRt7FX87YlwgH8w9kMENz/sqFAT7ex2Aw4FV1kuk5A+IkGKv6pUyDsyHAWnEFR
atAdZaRzPQ/oTTm6snx/LTgrcO5r/YEuKjQ8RII+qfB1Uj9wy2RvEMdLB92oic8+NV8NuS+Z0vja
MqIBQHL3oDxhvJVhq/bH5ZERgmSewEFyZDyG6NPanbRi2ol72yeXEpsnpaY+b7B/RS+nUbVQxdMh
qLJLnaBBT3MqBYnqbHwA6rTLY80Db6SQdp1INYWkWG/VSq1apJw2FU+E9SdtzEjIE5VhPtYL1iNX
42M0yU89SJD444E1eMPeye2pEcp7cVZy8jQsJFcppedEm9alR2I5z3I2QweNaj9G5E8CTfmv9yAQ
ju8FnFr73U9iQUTFntrP966B9byX7fK0bPIFeoAcyI6mvA+aTiGjR/Ru1S6ONOsY7CoUyvWMX6a1
fhXqL0oauM0HRbQoYBg/mKO24YqkI6KinLBYeWyiYVVY1aGFnUPt46aRJ3wmido5Um33JWCTzSrz
W0rhS9vsdo+AxC4TsDd4Wts+YiTDrOJiKHHis2c41RXTwKFbozRoOoFzuyMjEB+/5LDGSUECefxH
Xm7gCxyMrjAUPTeTUyRfRIgbqneYnSJPmu23pRXAnOk+SXnfb1E2XYXIXpsQrzcJwfoSp5l+hmb9
lTKYnvvo/aes9V9z6Wd0V8IbtfYlIJ7ZfgzU+ZM2ip6/FHlvUFbzqGeepZ4recJ2E39+YnW8FgCn
vHtZUyxO6PKyyHK2IPnkE8QrvBJ15j6Wp7AK/cTrDi0mZaktKuea+hPF0Ez+0vpVtYs6z7W/UiuI
n4BeuWfXUPJCE1Jow5ytZSTkNunVWQnw2yL48q6Wg2ybbdbuN257FRfTJanHJJjPfky3hrdtnccp
09s1QuFC2cFpgc38rkftrj+GemnO/FJ3MiXaMj9iaYwvZKUgguzmRP6Maw2I7wr8M9J87uPMwe4e
wr2kQEOwNDZG48psvRsk79i+CT6ZNahz57XjYHOlHJDHpvBl0aRT4QqhZfyaqeJFCWEbusalTrBm
TnfWzb7jjV1h7wefxeCyxk2DgfNqYTjrT+HemtfmvNnjMmahQIPXE0NRJNk7hI8aBNZU9b8z1nik
APfPCdrONAfBkY56Oy4V30iwyUhIMi057jffdS+chnmoZDqP4l3GP1+UINNLz9U7YVb4axL717dj
qx3ZGKniiu9Q32+NTJLsSOQYCFxh+IcOufBA4FPE+7VjzOtcx8c0tX4tkzB69k2oD/rBhhfWIpRk
8yAazW6KtSeRy1eP9jiifaRIYUH1tozPz3DC1L53OTdZeiPP+KR7Ck+zHwZrfcH19wjTL+ID7ihi
AvUiWEPNR52TQZvF/UQc66H5oopZoAliENtmQIrcgod+6Wjmx/e/xW5ytlo/f0hC6yXuJJA36x8g
NhAN7NDyL8gzlEBEggYidzfhlchRiCoUa7FbOuzNH4rj7yFi2/4xRGqY3bXrkECW4Uo2S4r5SzhJ
m20E7HxaIPOeZ2PaEu9udRXhJgiZVDHBcAkV0jzmKSdpxgTwKBK5+S2iAzSQuJsqgbE5NtCSeAvh
TkXMx2rlVBbaJ596zIMWEoM73nHvslml2hQQARt9y8KJTXUye2Ra+SnCaJ8Crd1GnzmV4gV3uRhq
4JPA9z5EaUFA1RBZTNK1Vr0pJpShcM7i9aRBvUmBYUjlXIL0xM1+uNu+TCb4EVnNqE6RjLzhC8fZ
R4BBfEwx0mBJOK7LSghCUlBFMg5B2lIjSRS0TeQR3XQWqsEmHuCprLDYXK9WTcvrrx7ViIBvtzEN
rxxQ0oQVf1EDlbS0agz/Tk+ccEWw2QFP5aXAc5hwPzrOGetyExbUBPeXx+zxs7PmFTP2PwQPVmMG
0WOli1cwW4GSM92zlJqKG628vEvhmssN6pV1oz8nrhmXTZSSzBC0s/pbxkEmfHAWec8KoIthPmf2
g1kAvRf4EpfW/nkt0T3Kqcx88RbeMsZaSyw8UEOjexFIjcGHtTIw0Ize+scm225ywyHArq6oqdM8
HePkJrLyZArOMCSdEUM3J0U85b8p8XmJICf1VPdggGXpEpvbb6e6wVrQ93lDS0lZO1vK80phHu7O
6G7+CrehcZCl8ESWP/j6a2tMwjLDXbpcpJe45Vid6TRDXXqwkZ5UCuPVJNy0oSCS0AuHLcfRCFBS
heNGGnW7FPcXXJd/t1W8808pCRkRMzse6IBfuXrjxQdstRh24KQgN5mWnLjTeErwNlg3/wJpj5uf
I8otaT9s2xhPISsKEEPvrzO843BYx8xBoL4WI8QVnl9Wa96qtaqAoEi0H0pjmjUWyK7sAzSjbe5L
br1MbSVs4vSvlNKVHj0u1XvfGljSN75rnGmOt+aM7tYZkaBCugamZtomZZfy+GO2hppKmJb21aAA
+YMHaqgK/sdQ2TmAXqi79oQ3lrjrZKPco8LfmNn6g9opNGLwsKeSJxZP3BoA9t+C+ANVYeHoN/Iw
DTLs0hHJpNbfBTRSk+jISJs6MRiLk0s6AJ/6ounnWwr3POwJd4FE15NqHtTp8uK+toAnVqMHrWz8
fFixyBv+H8ecqh+AwHQeB9uvJiP8JtQPteGzZcVt4PSf755iIT/bTlc5hudHP3Am96+BEqymWabp
22H/o1EXYGI3H0Pk/dtD8qqW8Pcvs9Dc/w5WD7ev3WqUdcIJj1Ju8az/04n7hLytjUKq9vAgUgEY
fXHa9yREAH52HR7aEsoG4u21BC4QweaO5WQB5fZd06q1xu3rYTO1QMilpg3dKHoI1HI7mqAEuyWl
pT6CIWCt4TRYL+1YnWqRPvc6FWqAD821/3eTJY1Kde8tvWRqx52GCWBPwFwGrhOwc6QINuMC5D+c
n7ll22rFK/Q+r8X0YYLS7sQ5kAQqNrTDXF02fnBwEemQ2aZHCcbOkVg7v9vy3HAhj5gX0pEGCuz3
Ntrv+W1nHEowYl0IC6r5y/WYP20fWkkO0n4zohyCFlDpJi11uB239Px3vkvgC3cbjFkcBJ5dnwM4
OytS3FDlNH5oLggvJ3Tk/V7tmQ2fZWLP2vgcaAYadoGZPJPoyPZM9oFn44aZj8q2kzrI23QiFpE2
j7tWN46WT/194Mvj2ql4RU7R+F2EumAG45LbELnwCKQv6jd8NQwWJcKtTNxdfypP9PsnOwGZ8qCY
iE4TY9abGzUg/S/EGMRzZdn+7uDpaeYWeAIVMu+wGszVOnWNst5Uv5tmH2sjLpaS3fthzzfKPdjR
dCr9wR/QFgc75DQqFZQf0jdktcNXJ4YE9Fn0k+GyBjjpCMO2G0yP/ISeaegPfqccEMgp9zB/sosL
JLf5XXoz9iW7HWw1OLu+OkB9lZ1wRODasdDcy4Ypc9xauswWaZD3PQawtehx4l6G+Zcd33muvFyH
2IwVK5FbYhV0GEtxdP3G7pw/noXM+W6aIk/xUVAxlWeZtUjTPr0gC27T/zaFeZ2SAKoex+s2vRF9
HsjbYIymeM/a1dWUVR9JVsFugBOSYV1lW4EkMVFR8VF/Anon4enw2b+ftBU6k2G2ta/3U3QLMVjM
S29TAKKJW1c2Mwu/b0uKzwnywtlB1LZ6tPaZrMZmxcXamorhrCQCPz0g5v2nEAqp9X896eIAQlMi
mUvTIDphOj1ffygz7wLtcVPckEbiAPnfjWxZLmV4IY16IfCmroZuNBv6UR5RiBssggu2sFO5Ti4e
cZ4+Y55Bcg3iUGJHCuOohOd0/KYBMZrpx+tjPKlE1eJGcRF6Kgp8EaBjZEMa0f5HnhkS1Tzl/y6Z
Tjk5jFHg/hmlXLKraojyqqlVV7S/uRG9VfGulThueLM+v+/EP4kUKijSUongdhKNZLyDIISRbAHF
CPXMTDa7u4KIiU1ywSbmANl4MZiNS/WetJ6BbQLUEIbkLccnBmZcFDoVZbSA6zuZXg8xoJOz7CUh
3QkPRe5YEoEouR9ZNl/hBa6TgmAIaHJJjd8FypjiMcff+CnH0/1VkNi0hWEF38FAmJaVPmxsuTx8
XEi+UYWeUNOuAZNYAOoPwMrlTP+ZID3rAXdReDZxvIyUdvhaL4LnNzbBGmy1r6u2O5IdaROWjoM7
1qKQswed/KVu8Ln2aW1PbFeb7MyPnlkoRxytkoUTDfI4ym9CfmqiNyNZVww9a55A0TIu9K7B9hSI
4zbvBGXp7rNOCfg/7yVdqEG0Ha0LUTBzsrx/oJ164lRZRUVGWbznVNLK9VEbVF1ko0YZXb/1hz0T
FqiSRC7hdFBYk0zudHnX+95y6kfwz2bYx0VoNrv5fokAqZcPP5wF5x09SakQD3aBPx/ig05Caacp
F+j4kJKsQ5MEwn7aTO51a2M3ftXjTeWDly3qvmt95VfNVt8sPC9vNepMCTTqRVxFy4kyJHRezmM+
4F6EV7GqJt5nurIvfxWmMiCofYBTDNLMeE/gC3SyommB5GxlhTS13Y1+IGcZBJxIxp9umSq0ICZO
eAOY6uceuufn1QQ5O0CjAnVr2FxVN+7WEQaA5JsQCatsZVI7D9I6OY+w3mPa1MsN8aaS4fAcaCLZ
56LkT+Ll/CDYAG83P8h22njGzx2LIaD+FEoOMydugYOAP2s5NyskzFL7xlRrc0Pge1bBKkmbKT7o
2iMfcd7p+eY75WrlxWRY4jm/LTZ2tII49/f2vCuKMGmBtKcKgILdmrf/JLQqRtsLje1iRLFpRkd+
usqw9UQQntyEpbUOIMfsPpx8AuEsQC75WuxoAb93fhIWkX3y5L9W5Y2ovTHQ+odQTLfuiG2tzNJn
3QqJp9yBTxsB+FU8gvy+CZ5FVhT4hoQKWulQNH7yAZiNHzldSnV3EKk+R5qXmJZbsv0zj8eUQudZ
5oVwdRsJ1CHGJ/OJ9hELkmJZgqleJEEr3SL7L/VvR43xJsTy8H7uCapNYPqvPdbeuABNaXlyTH42
cVhYrOZySUrY+EX9L4gASNzlZGwnVtXjAFAW5T2rxdPrN+nDivGcNCo1t6woLb8JsKgfsbk3DNCR
IL0cuDR6TRGnXCvvs68Qgi78VrLoQZcCI8wtkqsIY0ynY5sxP7jd1hzWB+k9u4Oqn54P0bWnWPC5
Pr1ZFF99rLoGChB3HSnAuZVUtzMsktyzgJsufd66dsBitp22SbcWiwArIpNgDYaIRcfA9ScsZVKj
ji8OdUlNwgmqHdarU1xChf16v6kphaTxFrnh5AWoKCOwdYhFJuLvcPDSOBFKuUMa7L33ljWtNkJ3
lsDkW3Kg1coDKIsnIpDGlN62NJkeKGcTGHK5TWKwnPbZBIMSga54OVr1ty3a2NUXdAfp2gGExgyS
qHZS1WOW8qbaxoNVXu/KSTAbx30Ue32cTNtqrR5G8yJUMQFOTgEpCQ3MD2zt531CnyWQf+XA+2nw
D1oPiXr9RY6Z+Qx8nycLrNTwZtyDnRF8BwykoFWjwK2olrzeZtzVrrSL7aVkEJeg24dzipqxtw3N
MtSEQhjx/oQdaY77A4fOqefa2Yh3IaJWLWa8tiDiY5cFjdjxZx9zOQZyRv8XsVUSwZxbpd4+3oaf
3fK8zcw2ipcq82KA+U8HT/rlnR6p0InOHBO5aMy5Mud5UqK/jkZqqtHVMiRbKRv9W0EWcnQmLo0h
IKFMx0we/nMxG7r86teBYqmcqe4nw5CWgHBNVSi8Nr/yEYVi06bnuFIKtKmyTuGwZ5AEGHoV181t
tBO/OOOA4VyMTb7VC75vXDTCpHSMqcUjQi0z8sKokG827Sg9Vj8nCLCpL1Z4moQcMjTdyiGrZc+z
CTdN3JuYfWOYCqViebrMEsh5f0W26IUzGvEO0gkjB7WbMRSiFeOUNm5iyXGA6+fXNnmdDJNz1hDV
mtA7eIXcJQm0SYZPo6WVhHVEoZLSOMjeLFgNzbDH1vDhyD1JLCfVvFo4DfZ+fhuFkbDEq5o7JEtN
pvwEU7NUeM3KLM7g1aEk3U6GahkGRD6Zupf3jJT8nsLuBnbQponqEmN86vTT5ySEFkUEIw89m8Wq
FsLjcK5WCbZC2bGrM9kHpJ9jK6PIuAZJqHyWjiuaSQd+YcZc89ZmXnMquEWOWepsKdsosNIlpS9L
Sk76a/qU5z/fmuNP8f/8fkh9C92i2VfxDrzJbJcRjEcuUMLnt9cratfp+WykBciPj8+VCQa/AJTX
Jn5nfNAwtbPaZVzwaDoCj4VcqkTob6w2KtiOrQ==
`protect end_protected
